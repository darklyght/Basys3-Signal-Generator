`timescale 1ns / 1ps

module character_rom(
    input CLK,
    input CHANNEL,
    input DC,
    input MIN_MAX,
    input BOTH,
    input WAVE,
    input AMP_MODE,
    input [39:0] FREQ1,
    input [31:0] MAX_AMP1,
    input [31:0] MIN_AMP1,
    input [1:0] WAVE1,
    input [1:0] FORM1,
    input [39:0] FREQ2,
    input [31:0] MAX_AMP2,
    input [31:0] MIN_AMP2,
    input [1:0] WAVE2,
    input [1:0] FORM2,
    input KEYBOARD,
    input MAX_AMP_MOD,
    input MIN_MAX_AMP_MOD,
    input FREQ_MOD,
    input [23:0] BANDWIDTH,
    input PHASE_MOD,
    input [23:0] DUTY_CYCLE,
    input SUPERPOSE,
    input [4:0] ROW,
    input [6:0] COL,
    output reg [7:0] DATA
    );
    
    reg [4:0] ROW_REG;
    reg [6:0] COL_REG;
    
    always @ (posedge CLK) begin
        ROW_REG <= ROW;
        COL_REG <= COL;
    end
    
    always @ (*) begin
        case ({ROW_REG, COL_REG})
            // Row 0
            12'b00000_0000000: DATA = 8'h44;
            12'b00000_0000001: DATA = 8'h41;
            12'b00000_0000010: DATA = 8'h52;
            12'b00000_0000011: DATA = 8'h4B;
            12'b00000_0000100: DATA = 8'h4C;
            12'b00000_0000101: DATA = 8'h59;
            12'b00000_0000110: DATA = 8'h47;
            12'b00000_0000111: DATA = 8'h48;
            12'b00000_0001000: DATA = 8'h54;
            12'b00000_0001001: DATA = 8'h27;
            12'b00000_0001010: DATA = 8'h53;
            12'b00000_0001011: DATA = 8'h00;
            12'b00000_0001100: DATA = 8'h53;
            12'b00000_0001101: DATA = 8'h49;
            12'b00000_0001110: DATA = 8'h47;
            12'b00000_0001111: DATA = 8'h4E;
            12'b00000_0010000: DATA = 8'h41;
            12'b00000_0010001: DATA = 8'h4C;
            12'b00000_0010010: DATA = 8'h00;
            12'b00000_0010011: DATA = 8'h47;
            12'b00000_0010100: DATA = 8'h45;
            12'b00000_0010101: DATA = 8'h4E;
            12'b00000_0010110: DATA = 8'h45;
            12'b00000_0010111: DATA = 8'h52;
            12'b00000_0011000: DATA = 8'h41;
            12'b00000_0011001: DATA = 8'h54;
            12'b00000_0011010: DATA = 8'h4F;
            12'b00000_0011011: DATA = 8'h52;
            12'b00000_0011100: DATA = 8'h00;
            12'b00000_0011101: DATA = 8'h00;
            12'b00000_0011110: DATA = 8'h00;
            12'b00000_0011111: DATA = 8'h00;
            12'b00000_0100000: DATA = 8'h00;
            12'b00000_0100001: DATA = 8'h00;
            12'b00000_0100010: DATA = 8'h00;
            12'b00000_0100011: DATA = 8'h00;
            12'b00000_0100100: DATA = 8'h00;
            12'b00000_0100101: DATA = 8'h00;
            12'b00000_0100110: DATA = 8'h00;
            12'b00000_0100111: DATA = 8'h00;
            12'b00000_0101000: DATA = 8'h00;
            12'b00000_0101001: DATA = 8'h00;
            12'b00000_0101010: DATA = 8'h00;
            12'b00000_0101011: DATA = 8'h00;
            12'b00000_0101100: DATA = 8'h00;
            12'b00000_0101101: DATA = 8'h00;
            12'b00000_0101110: DATA = 8'h00;
            12'b00000_0101111: DATA = 8'h00;
            12'b00000_0110000: DATA = 8'h00;
            12'b00000_0110001: DATA = 8'h00;
            12'b00000_0110010: DATA = 8'h00;
            12'b00000_0110011: DATA = 8'h00;
            12'b00000_0110100: DATA = 8'h00;
            12'b00000_0110101: DATA = 8'h00;
            12'b00000_0110110: DATA = 8'h00;
            12'b00000_0110111: DATA = 8'h00;
            12'b00000_0111000: DATA = 8'h00;
            12'b00000_0111001: DATA = 8'h00;
            12'b00000_0111010: DATA = 8'h00;
            12'b00000_0111011: DATA = 8'h00;
            12'b00000_0111100: DATA = 8'h00;
            12'b00000_0111101: DATA = 8'h00;
            12'b00000_0111110: DATA = 8'h00;
            12'b00000_0111111: DATA = 8'h00;
            12'b00000_1000000: DATA = 8'h00;
            12'b00000_1000001: DATA = 8'h00;
            12'b00000_1000010: DATA = 8'h00;
            12'b00000_1000011: DATA = 8'h00;
            12'b00000_1000100: DATA = 8'h00;
            12'b00000_1000101: DATA = 8'h00;
            12'b00000_1000110: DATA = 8'h00;
            12'b00000_1000111: DATA = 8'h00;
            12'b00000_1001000: DATA = 8'h00;
            12'b00000_1001001: DATA = 8'h00;
            12'b00000_1001010: DATA = 8'h00;
            12'b00000_1001011: DATA = 8'h00;
            12'b00000_1001100: DATA = 8'h00;
            12'b00000_1001101: DATA = 8'h00;
            12'b00000_1001110: DATA = 8'h00;
            12'b00000_1001111: DATA = 8'h00;
            // Row 1
            12'b00001_0000000: DATA = 8'h00;
            12'b00001_0000001: DATA = 8'h00;
            12'b00001_0000010: DATA = 8'h00;
            12'b00001_0000011: DATA = 8'h00;
            12'b00001_0000100: DATA = 8'h00;
            12'b00001_0000101: DATA = 8'h00;
            12'b00001_0000110: DATA = 8'h00;
            12'b00001_0000111: DATA = 8'h00;
            12'b00001_0001000: DATA = 8'h00;
            12'b00001_0001001: DATA = 8'h00;
            12'b00001_0001010: DATA = 8'h00;
            12'b00001_0001011: DATA = 8'h00;
            12'b00001_0001100: DATA = 8'h00;
            12'b00001_0001101: DATA = 8'h00;
            12'b00001_0001110: DATA = 8'h00;
            12'b00001_0001111: DATA = 8'h00;
            12'b00001_0010000: DATA = 8'h00;
            12'b00001_0010001: DATA = 8'h00;
            12'b00001_0010010: DATA = 8'h00;
            12'b00001_0010011: DATA = 8'h00;
            12'b00001_0010100: DATA = 8'h00;
            12'b00001_0010101: DATA = 8'h00;
            12'b00001_0010110: DATA = 8'h00;
            12'b00001_0010111: DATA = 8'h00;
            12'b00001_0011000: DATA = 8'h00;
            12'b00001_0011001: DATA = 8'h00;
            12'b00001_0011010: DATA = 8'h00;
            12'b00001_0011011: DATA = 8'h00;
            12'b00001_0011100: DATA = 8'h00;
            12'b00001_0011101: DATA = 8'h00;
            12'b00001_0011110: DATA = 8'h00;
            12'b00001_0011111: DATA = 8'h00;
            12'b00001_0100000: DATA = 8'h00;
            12'b00001_0100001: DATA = 8'h00;
            12'b00001_0100010: DATA = 8'h00;
            12'b00001_0100011: DATA = 8'h00;
            12'b00001_0100100: DATA = 8'h00;
            12'b00001_0100101: DATA = 8'h00;
            12'b00001_0100110: DATA = 8'h00;
            12'b00001_0100111: DATA = 8'h00;
            12'b00001_0101000: DATA = 8'h00;
            12'b00001_0101001: DATA = 8'h00;
            12'b00001_0101010: DATA = 8'h00;
            12'b00001_0101011: DATA = 8'h00;
            12'b00001_0101100: DATA = 8'h00;
            12'b00001_0101101: DATA = 8'h00;
            12'b00001_0101110: DATA = 8'h00;
            12'b00001_0101111: DATA = 8'h00;
            12'b00001_0110000: DATA = 8'h00;
            12'b00001_0110001: DATA = 8'h00;
            12'b00001_0110010: DATA = 8'h00;
            12'b00001_0110011: DATA = 8'h00;
            12'b00001_0110100: DATA = 8'h00;
            12'b00001_0110101: DATA = 8'h00;
            12'b00001_0110110: DATA = 8'h00;
            12'b00001_0110111: DATA = 8'h00;
            12'b00001_0111000: DATA = 8'h00;
            12'b00001_0111001: DATA = 8'h00;
            12'b00001_0111010: DATA = 8'h00;
            12'b00001_0111011: DATA = 8'h00;
            12'b00001_0111100: DATA = 8'h00;
            12'b00001_0111101: DATA = 8'h00;
            12'b00001_0111110: DATA = 8'h00;
            12'b00001_0111111: DATA = 8'h00;
            12'b00001_1000000: DATA = 8'h00;
            12'b00001_1000001: DATA = 8'h00;
            12'b00001_1000010: DATA = 8'h00;
            12'b00001_1000011: DATA = 8'h00;
            12'b00001_1000100: DATA = 8'h00;
            12'b00001_1000101: DATA = 8'h00;
            12'b00001_1000110: DATA = 8'h00;
            12'b00001_1000111: DATA = 8'h00;
            12'b00001_1001000: DATA = 8'h00;
            12'b00001_1001001: DATA = 8'h00;
            12'b00001_1001010: DATA = 8'h00;
            12'b00001_1001011: DATA = 8'h00;
            12'b00001_1001100: DATA = 8'h00;
            12'b00001_1001101: DATA = 8'h00;
            12'b00001_1001110: DATA = 8'h00;
            12'b00001_1001111: DATA = 8'h00;
            // Row 2
            12'b00010_0000000: DATA = 8'h43;
            12'b00010_0000001: DATA = 8'h48;
            12'b00010_0000010: DATA = 8'h41;
            12'b00010_0000011: DATA = 8'h4E;
            12'b00010_0000100: DATA = 8'h4E;
            12'b00010_0000101: DATA = 8'h45;
            12'b00010_0000110: DATA = 8'h4C;
            12'b00010_0000111: DATA = 8'h00;
            12'b00010_0001000: DATA = 8'h31;
            12'b00010_0001001: DATA = 8'h00;
            12'b00010_0001010: DATA = (CHANNEL == 0) ? 8'h3C : 8'h00;
            12'b00010_0001011: DATA = 8'h00;
            12'b00010_0001100: DATA = (CHANNEL == 0 && DC == 1) ? 8'h44 : 8'h00;
            12'b00010_0001101: DATA = (CHANNEL == 0 && DC == 1) ? 8'h43 : 8'h00;
            12'b00010_0001110: DATA = 8'h00;
            12'b00010_0001111: DATA = 8'h00;
            12'b00010_0010000: DATA = 8'h00;
            12'b00010_0010001: DATA = 8'h00;
            12'b00010_0010010: DATA = 8'h00;
            12'b00010_0010011: DATA = 8'h00;
            12'b00010_0010100: DATA = 8'h00;
            12'b00010_0010101: DATA = 8'h00;
            12'b00010_0010110: DATA = 8'h00;
            12'b00010_0010111: DATA = 8'h00;
            12'b00010_0011000: DATA = 8'h00;
            12'b00010_0011001: DATA = 8'h00;
            12'b00010_0011010: DATA = 8'h00;
            12'b00010_0011011: DATA = 8'h00;
            12'b00010_0011100: DATA = 8'hD4;
            12'b00010_0011101: DATA = 8'hC8;
            12'b00010_0011110: DATA = 8'hC8;
            12'b00010_0011111: DATA = 8'hC8;
            12'b00010_0100000: DATA = 8'hC8;
            12'b00010_0100001: DATA = 8'hC8;
            12'b00010_0100010: DATA = 8'hC8;
            12'b00010_0100011: DATA = 8'hC8;
            12'b00010_0100100: DATA = 8'hC8;
            12'b00010_0100101: DATA = 8'hC8;
            12'b00010_0100110: DATA = 8'hC8;
            12'b00010_0100111: DATA = 8'hD5;
            12'b00010_0101000: DATA = 8'h00;
            12'b00010_0101001: DATA = 8'h00;
            12'b00010_0101010: DATA = 8'h00;
            12'b00010_0101011: DATA = 8'h00;
            12'b00010_0101100: DATA = 8'h00;
            12'b00010_0101101: DATA = 8'h00;
            12'b00010_0101110: DATA = 8'h00;
            12'b00010_0101111: DATA = 8'h00;
            12'b00010_0110000: DATA = 8'h00;
            12'b00010_0110001: DATA = 8'h00;
            12'b00010_0110010: DATA = 8'h00;
            12'b00010_0110011: DATA = 8'h00;
            12'b00010_0110100: DATA = 8'h00;
            12'b00010_0110101: DATA = 8'h00;
            12'b00010_0110110: DATA = 8'h00;
            12'b00010_0110111: DATA = 8'h00;
            12'b00010_0111000: DATA = 8'h00;
            12'b00010_0111001: DATA = 8'h00;
            12'b00010_0111010: DATA = 8'h00;
            12'b00010_0111011: DATA = 8'h00;
            12'b00010_0111100: DATA = 8'h00;
            12'b00010_0111101: DATA = 8'h00;
            12'b00010_0111110: DATA = 8'h00;
            12'b00010_0111111: DATA = 8'h00;
            12'b00010_1000000: DATA = 8'h00;
            12'b00010_1000001: DATA = 8'h00;
            12'b00010_1000010: DATA = 8'h00;
            12'b00010_1000011: DATA = 8'h00;
            12'b00010_1000100: DATA = 8'h00;
            12'b00010_1000101: DATA = 8'h00;
            12'b00010_1000110: DATA = 8'h00;
            12'b00010_1000111: DATA = 8'h00;
            12'b00010_1001000: DATA = 8'h00;
            12'b00010_1001001: DATA = 8'h00;
            12'b00010_1001010: DATA = 8'h00;
            12'b00010_1001011: DATA = 8'h00;
            12'b00010_1001100: DATA = 8'h00;
            12'b00010_1001101: DATA = 8'h00;
            12'b00010_1001110: DATA = 8'h00;
            12'b00010_1001111: DATA = 8'h00;
            // Row 3
            12'b00011_0000000: DATA = 8'h46;
            12'b00011_0000001: DATA = 8'h52;
            12'b00011_0000010: DATA = 8'h45;
            12'b00011_0000011: DATA = 8'h51;
            12'b00011_0000100: DATA = 8'h55;
            12'b00011_0000101: DATA = 8'h45;
            12'b00011_0000110: DATA = 8'h4E;
            12'b00011_0000111: DATA = 8'h43;
            12'b00011_0001000: DATA = 8'h59;
            12'b00011_0001001: DATA = 8'h00;
            12'b00011_0001010: DATA = 8'h00;
            12'b00011_0001011: DATA = 8'h00;
            12'b00011_0001100: DATA = 8'h00;
            12'b00011_0001101: DATA = 8'h00;
            12'b00011_0001110: DATA = FREQ1[39:32];
            12'b00011_0001111: DATA = FREQ1[31:24];
            12'b00011_0010000: DATA = FREQ1[23:16];
            12'b00011_0010001: DATA = FREQ1[15:8];
            12'b00011_0010010: DATA = FREQ1[7:0];
            12'b00011_0010011: DATA = 8'h00;
            12'b00011_0010100: DATA = 8'h00;
            12'b00011_0010101: DATA = 8'h00;
            12'b00011_0010110: DATA = 8'h00;
            12'b00011_0010111: DATA = 8'h00;
            12'b00011_0011000: DATA = 8'h00;
            12'b00011_0011001: DATA = 8'h00;
            12'b00011_0011010: DATA = 8'h00;
            12'b00011_0011011: DATA = 8'h00;
            12'b00011_0011100: DATA = 8'hC6;
            12'b00011_0011101: DATA = (FORM1 == 2'b10) ? 8'h00 : (WAVE1 == 2'b00) ? 8'h94 : (WAVE1 == 2'b01) ? 8'hBC : (WAVE1 == 2'b10) ? 8'hA8 : 8'h80;
            12'b00011_0011110: DATA = (FORM1 == 2'b10) ? 8'h00 : (WAVE1 == 2'b00) ? 8'h95 : (WAVE1 == 2'b01) ? 8'hBD : (WAVE1 == 2'b10) ? 8'hA9 : 8'h81;
            12'b00011_0011111: DATA = (FORM1 == 2'b10) ? 8'h00 : (WAVE1 == 2'b00) ? 8'h96 : (WAVE1 == 2'b01) ? 8'hBE : (WAVE1 == 2'b10) ? 8'hAA : 8'h82;
            12'b00011_0100000: DATA = (FORM1 == 2'b10) ? 8'h00 : (WAVE1 == 2'b00) ? 8'h97 : (WAVE1 == 2'b01) ? 8'hBF : (WAVE1 == 2'b10) ? 8'hAB : 8'h83;
            12'b00011_0100001: DATA = (FORM1 == 2'b10) ? 8'h00 : (WAVE1 == 2'b00) ? 8'h98 : (WAVE1 == 2'b01) ? 8'hC0 : (WAVE1 == 2'b10) ? 8'hAC : 8'h84;
            12'b00011_0100010: DATA = (FORM1 == 2'b00) ? 8'h00 : (FORM1 == 2'b01) ? 8'h00 : (WAVE1 == 2'b00) ? 8'h94 : (WAVE1 == 2'b01) ? 8'hD8 : (WAVE1 == 2'b10) ? 8'hA8 : 8'h80;
            12'b00011_0100011: DATA = (FORM1 == 2'b00) ? 8'h00 : (FORM1 == 2'b01) ? 8'h00 : (WAVE1 == 2'b00) ? 8'h95 : (WAVE1 == 2'b01) ? 8'hD9 : (WAVE1 == 2'b10) ? 8'hA9 : 8'h81;
            12'b00011_0100100: DATA = (FORM1 == 2'b00) ? 8'h00 : (FORM1 == 2'b01) ? 8'h00 : (WAVE1 == 2'b00) ? 8'h96 : (WAVE1 == 2'b01) ? 8'hDA : (WAVE1 == 2'b10) ? 8'hAA : 8'h82;
            12'b00011_0100101: DATA = (FORM1 == 2'b00) ? 8'h00 : (FORM1 == 2'b01) ? 8'h00 : (WAVE1 == 2'b00) ? 8'h97 : (WAVE1 == 2'b01) ? 8'hDB : (WAVE1 == 2'b10) ? 8'hAB : 8'h83;
            12'b00011_0100110: DATA = (FORM1 == 2'b00) ? 8'h00 : (FORM1 == 2'b01) ? 8'h00 : (WAVE1 == 2'b00) ? 8'h98 : (WAVE1 == 2'b01) ? 8'hDC : (WAVE1 == 2'b10) ? 8'hAC : 8'h84;
            12'b00011_0100111: DATA = 8'hC7;
            12'b00011_0101000: DATA = 8'h00;
            12'b00011_0101001: DATA = 8'h00;
            12'b00011_0101010: DATA = 8'h00;
            12'b00011_0101011: DATA = 8'h00;
            12'b00011_0101100: DATA = 8'h00;
            12'b00011_0101101: DATA = 8'h00;
            12'b00011_0101110: DATA = 8'h00;
            12'b00011_0101111: DATA = 8'h00;
            12'b00011_0110000: DATA = 8'h00;
            12'b00011_0110001: DATA = 8'h00;
            12'b00011_0110010: DATA = 8'h00;
            12'b00011_0110011: DATA = 8'h00;
            12'b00011_0110100: DATA = 8'h00;
            12'b00011_0110101: DATA = 8'h00;
            12'b00011_0110110: DATA = 8'h00;
            12'b00011_0110111: DATA = 8'h00;
            12'b00011_0111000: DATA = 8'h00;
            12'b00011_0111001: DATA = 8'h00;
            12'b00011_0111010: DATA = 8'h00;
            12'b00011_0111011: DATA = 8'h00;
            12'b00011_0111100: DATA = 8'h00;
            12'b00011_0111101: DATA = 8'h00;
            12'b00011_0111110: DATA = 8'h00;
            12'b00011_0111111: DATA = 8'h00;
            12'b00011_1000000: DATA = 8'h00;
            12'b00011_1000001: DATA = 8'h00;
            12'b00011_1000010: DATA = 8'h00;
            12'b00011_1000011: DATA = 8'h00;
            12'b00011_1000100: DATA = 8'h00;
            12'b00011_1000101: DATA = 8'h00;
            12'b00011_1000110: DATA = 8'h00;
            12'b00011_1000111: DATA = 8'h00;
            12'b00011_1001000: DATA = 8'h00;
            12'b00011_1001001: DATA = 8'h00;
            12'b00011_1001010: DATA = 8'h00;
            12'b00011_1001011: DATA = 8'h00;
            12'b00011_1001100: DATA = 8'h00;
            12'b00011_1001101: DATA = 8'h00;
            12'b00011_1001110: DATA = 8'h00;
            12'b00011_1001111: DATA = 8'h00;
            // Row 4
            12'b00100_0000000: DATA = 8'h4D;
            12'b00100_0000001: DATA = 8'h41;
            12'b00100_0000010: DATA = 8'h58;
            12'b00100_0000011: DATA = 8'h00;
            12'b00100_0000100: DATA = 8'h41;
            12'b00100_0000101: DATA = 8'h4D;
            12'b00100_0000110: DATA = 8'h50;
            12'b00100_0000111: DATA = 8'h4C;
            12'b00100_0001000: DATA = 8'h49;
            12'b00100_0001001: DATA = 8'h54;
            12'b00100_0001010: DATA = 8'h55;
            12'b00100_0001011: DATA = 8'h44;
            12'b00100_0001100: DATA = 8'h45;
            12'b00100_0001101: DATA = 8'h00;
            12'b00100_0001110: DATA = MAX_AMP1[31:24];
            12'b00100_0001111: DATA = (AMP_MODE == 1) ? MAX_AMP1[23:16] : 8'h2E;
            12'b00100_0010000: DATA = (AMP_MODE == 1) ? MAX_AMP1[15:8] : MAX_AMP1[23:16];
            12'b00100_0010001: DATA = (AMP_MODE == 1) ? MAX_AMP1[7:0] : MAX_AMP1[15:8];
            12'b00100_0010010: DATA = (AMP_MODE == 1) ? 8'h00 : MAX_AMP1[7:0];
            12'b00100_0010011: DATA = 8'h00;
            12'b00100_0010100: DATA = 8'h00;
            12'b00100_0010101: DATA = 8'h00;
            12'b00100_0010110: DATA = 8'h00;
            12'b00100_0010111: DATA = 8'h00;
            12'b00100_0011000: DATA = 8'h00;
            12'b00100_0011001: DATA = 8'h00;
            12'b00100_0011010: DATA = 8'h00;
            12'b00100_0011011: DATA = 8'h00;
            12'b00100_0011100: DATA = 8'hC6;
            12'b00100_0011101: DATA = (FORM1 == 2'b10) ? 8'h00 : (WAVE1 == 2'b00) ? 8'h99 : (WAVE1 == 2'b01) ? 8'hC1 : (WAVE1 == 2'b10) ? 8'hAD : 8'h85;
            12'b00100_0011110: DATA = (FORM1 == 2'b10) ? 8'h00 : (WAVE1 == 2'b00) ? 8'h9A : (WAVE1 == 2'b01) ? 8'hC2 : (WAVE1 == 2'b10) ? 8'hAE : 8'h86;
            12'b00100_0011111: DATA = (FORM1 == 2'b10) ? 8'h00 : (WAVE1 == 2'b00) ? 8'h9B : (WAVE1 == 2'b01) ? 8'hC3 : (WAVE1 == 2'b10) ? 8'hAF : 8'h87;
            12'b00100_0100000: DATA = (FORM1 == 2'b10) ? 8'h00 : (WAVE1 == 2'b00) ? 8'h9C : (WAVE1 == 2'b01) ? 8'hC4 : (WAVE1 == 2'b10) ? 8'hB0 : 8'h88;
            12'b00100_0100001: DATA = (FORM1 == 2'b10) ? 8'h00 : (WAVE1 == 2'b00) ? 8'h9D : (WAVE1 == 2'b01) ? 8'hC5 : (WAVE1 == 2'b10) ? 8'hB1 : 8'h89;
            12'b00100_0100010: DATA = (FORM1 == 2'b00) ? 8'h00 : (FORM1 == 2'b01) ? 8'h00 : (WAVE1 == 2'b00) ? 8'h99 : (WAVE1 == 2'b01) ? 8'hDD : (WAVE1 == 2'b10) ? 8'hAD : 8'h85;
            12'b00100_0100011: DATA = (FORM1 == 2'b00) ? 8'h00 : (FORM1 == 2'b01) ? 8'h00 : (WAVE1 == 2'b00) ? 8'h9A : (WAVE1 == 2'b01) ? 8'hDE : (WAVE1 == 2'b10) ? 8'hAE : 8'h86;
            12'b00100_0100100: DATA = (FORM1 == 2'b00) ? 8'h00 : (FORM1 == 2'b01) ? 8'h00 : (WAVE1 == 2'b00) ? 8'h9B : (WAVE1 == 2'b01) ? 8'hDF : (WAVE1 == 2'b10) ? 8'hAF : 8'h87;
            12'b00100_0100101: DATA = (FORM1 == 2'b00) ? 8'h00 : (FORM1 == 2'b01) ? 8'h00 : (WAVE1 == 2'b00) ? 8'h9C : (WAVE1 == 2'b01) ? 8'hE0 : (WAVE1 == 2'b10) ? 8'hB0 : 8'h88;
            12'b00100_0100110: DATA = (FORM1 == 2'b00) ? 8'h00 : (FORM1 == 2'b01) ? 8'h00 : (WAVE1 == 2'b00) ? 8'h9D : (WAVE1 == 2'b01) ? 8'hE1 : (WAVE1 == 2'b10) ? 8'hB1 : 8'h89;
            12'b00100_0100111: DATA = 8'hC7;
            12'b00100_0101000: DATA = 8'h00;
            12'b00100_0101001: DATA = 8'h00;
            12'b00100_0101010: DATA = 8'h00;
            12'b00100_0101011: DATA = 8'h00;
            12'b00100_0101100: DATA = 8'h00;
            12'b00100_0101101: DATA = 8'h00;
            12'b00100_0101110: DATA = 8'h00;
            12'b00100_0101111: DATA = 8'h00;
            12'b00100_0110000: DATA = 8'h00;
            12'b00100_0110001: DATA = 8'h00;
            12'b00100_0110010: DATA = 8'h00;
            12'b00100_0110011: DATA = 8'h00;
            12'b00100_0110100: DATA = 8'h00;
            12'b00100_0110101: DATA = 8'h00;
            12'b00100_0110110: DATA = 8'h00;
            12'b00100_0110111: DATA = 8'h00;
            12'b00100_0111000: DATA = 8'h00;
            12'b00100_0111001: DATA = 8'h00;
            12'b00100_0111010: DATA = 8'h00;
            12'b00100_0111011: DATA = 8'h00;
            12'b00100_0111100: DATA = 8'h00;
            12'b00100_0111101: DATA = 8'h00;
            12'b00100_0111110: DATA = 8'h00;
            12'b00100_0111111: DATA = 8'h00;
            12'b00100_1000000: DATA = 8'h00;
            12'b00100_1000001: DATA = 8'h00;
            12'b00100_1000010: DATA = 8'h00;
            12'b00100_1000011: DATA = 8'h00;
            12'b00100_1000100: DATA = 8'h00;
            12'b00100_1000101: DATA = 8'h00;
            12'b00100_1000110: DATA = 8'h00;
            12'b00100_1000111: DATA = 8'h00;
            12'b00100_1001000: DATA = 8'h00;
            12'b00100_1001001: DATA = 8'h00;
            12'b00100_1001010: DATA = 8'h00;
            12'b00100_1001011: DATA = 8'h00;
            12'b00100_1001100: DATA = 8'h00;
            12'b00100_1001101: DATA = 8'h00;
            12'b00100_1001110: DATA = 8'h00;
            12'b00100_1001111: DATA = 8'h00;
            // Row 5
            12'b00101_0000000: DATA = 8'h4D;
            12'b00101_0000001: DATA = 8'h49;
            12'b00101_0000010: DATA = 8'h4E;
            12'b00101_0000011: DATA = 8'h00;
            12'b00101_0000100: DATA = 8'h41;
            12'b00101_0000101: DATA = 8'h4D;
            12'b00101_0000110: DATA = 8'h50;
            12'b00101_0000111: DATA = 8'h4C;
            12'b00101_0001000: DATA = 8'h49;
            12'b00101_0001001: DATA = 8'h54;
            12'b00101_0001010: DATA = 8'h55;
            12'b00101_0001011: DATA = 8'h44;
            12'b00101_0001100: DATA = 8'h45;
            12'b00101_0001101: DATA = 8'h00;
            12'b00101_0001110: DATA = MIN_AMP1[31:24];
            12'b00101_0001111: DATA = (AMP_MODE == 1) ? MIN_AMP1[23:16] : 8'h2E;
            12'b00101_0010000: DATA = (AMP_MODE == 1) ? MIN_AMP1[15:8] : MIN_AMP1[23:16];
            12'b00101_0010001: DATA = (AMP_MODE == 1) ? MIN_AMP1[7:0] : MIN_AMP1[15:8];
            12'b00101_0010010: DATA = (AMP_MODE == 1) ? 8'h00 : MIN_AMP1[7:0];
            12'b00101_0010011: DATA = 8'h00;
            12'b00101_0010100: DATA = 8'h00;
            12'b00101_0010101: DATA = 8'h00;
            12'b00101_0010110: DATA = 8'h00;
            12'b00101_0010111: DATA = 8'h00;
            12'b00101_0011000: DATA = 8'h00;
            12'b00101_0011001: DATA = 8'h00;
            12'b00101_0011010: DATA = 8'h00;
            12'b00101_0011011: DATA = 8'h00;
            12'b00101_0011100: DATA = 8'hC6;
            12'b00101_0011101: DATA = (FORM1 == 2'b10 && WAVE1 == 2'b00) ? 8'h9E : (FORM1 == 2'b10 && WAVE1 == 2'b01) ? 8'hE2 : (FORM1 == 2'b10 && WAVE1 == 2'b10) ? 8'hB2 : (FORM1 == 2'b10 && WAVE1 == 2'b11) ? 8'h8A : 8'h00;
            12'b00101_0011110: DATA = (FORM1 == 2'b10 && WAVE1 == 2'b00) ? 8'h9F : (FORM1 == 2'b10 && WAVE1 == 2'b01) ? 8'hE3 : (FORM1 == 2'b10 && WAVE1 == 2'b10) ? 8'hB3 : (FORM1 == 2'b10 && WAVE1 == 2'b11) ? 8'h8B : 8'h00;
            12'b00101_0011111: DATA = (FORM1 == 2'b10 && WAVE1 == 2'b00) ? 8'hA0 : (FORM1 == 2'b10 && WAVE1 == 2'b01) ? 8'hE4 : (FORM1 == 2'b10 && WAVE1 == 2'b10) ? 8'hB4 : (FORM1 == 2'b10 && WAVE1 == 2'b11) ? 8'h8C : 8'h00;
            12'b00101_0100000: DATA = (FORM1 == 2'b10 && WAVE1 == 2'b00) ? 8'hA1 : (FORM1 == 2'b10 && WAVE1 == 2'b01) ? 8'hE5 : (FORM1 == 2'b10 && WAVE1 == 2'b10) ? 8'hB5 : (FORM1 == 2'b10 && WAVE1 == 2'b11) ? 8'h8D : 8'h00;
            12'b00101_0100001: DATA = (FORM1 == 2'b10 && WAVE1 == 2'b00) ? 8'hA2 : (FORM1 == 2'b10 && WAVE1 == 2'b01) ? 8'hE6 : (FORM1 == 2'b10 && WAVE1 == 2'b10) ? 8'hB6 : (FORM1 == 2'b10 && WAVE1 == 2'b11) ? 8'h8E : 8'h00;
            12'b00101_0100010: DATA = (FORM1 == 2'b01) ? 8'hC8 : (FORM1 == 2'b00 && WAVE1 == 2'b00) ? 8'h9E : (FORM1 == 2'b00 && WAVE1 == 2'b01) ? 8'hCA : (FORM1 == 2'b00 && WAVE1 == 2'b10) ? 8'hB2 : (FORM1 == 2'b00 && WAVE1 == 2'b11) ? 8'h8A : 8'h00;
            12'b00101_0100011: DATA = (FORM1 == 2'b01) ? 8'hC8 : (FORM1 == 2'b00 && WAVE1 == 2'b00) ? 8'h9F : (FORM1 == 2'b00 && WAVE1 == 2'b01) ? 8'hCB : (FORM1 == 2'b00 && WAVE1 == 2'b10) ? 8'hB3 : (FORM1 == 2'b00 && WAVE1 == 2'b11) ? 8'h8B : 8'h00;
            12'b00101_0100100: DATA = (FORM1 == 2'b01) ? 8'hC8 : (FORM1 == 2'b00 && WAVE1 == 2'b00) ? 8'hA0 : (FORM1 == 2'b00 && WAVE1 == 2'b01) ? 8'hCC : (FORM1 == 2'b00 && WAVE1 == 2'b10) ? 8'hB4 : (FORM1 == 2'b00 && WAVE1 == 2'b11) ? 8'h8C : 8'h00;
            12'b00101_0100101: DATA = (FORM1 == 2'b01) ? 8'hC8 : (FORM1 == 2'b00 && WAVE1 == 2'b00) ? 8'hA1 : (FORM1 == 2'b00 && WAVE1 == 2'b01) ? 8'hCD : (FORM1 == 2'b00 && WAVE1 == 2'b10) ? 8'hB5 : (FORM1 == 2'b00 && WAVE1 == 2'b11) ? 8'h8D : 8'h00;
            12'b00101_0100110: DATA = (FORM1 == 2'b01) ? 8'hC8 : (FORM1 == 2'b00 && WAVE1 == 2'b00) ? 8'hA2 : (FORM1 == 2'b00 && WAVE1 == 2'b01) ? 8'hCE : (FORM1 == 2'b00 && WAVE1 == 2'b10) ? 8'hB6 : (FORM1 == 2'b00 && WAVE1 == 2'b11) ? 8'h8E : 8'h00;
            12'b00101_0100111: DATA = 8'hC7;
            12'b00101_0101000: DATA = 8'h00;
            12'b00101_0101001: DATA = 8'h00;
            12'b00101_0101010: DATA = 8'h00;
            12'b00101_0101011: DATA = 8'h00;
            12'b00101_0101100: DATA = 8'h00;
            12'b00101_0101101: DATA = 8'h00;
            12'b00101_0101110: DATA = 8'h00;
            12'b00101_0101111: DATA = 8'h00;
            12'b00101_0110000: DATA = 8'h00;
            12'b00101_0110001: DATA = 8'h00;
            12'b00101_0110010: DATA = 8'h00;
            12'b00101_0110011: DATA = 8'h00;
            12'b00101_0110100: DATA = 8'h00;
            12'b00101_0110101: DATA = 8'h00;
            12'b00101_0110110: DATA = 8'h00;
            12'b00101_0110111: DATA = 8'h00;
            12'b00101_0111000: DATA = 8'h00;
            12'b00101_0111001: DATA = 8'h00;
            12'b00101_0111010: DATA = 8'h00;
            12'b00101_0111011: DATA = 8'h00;
            12'b00101_0111100: DATA = 8'h00;
            12'b00101_0111101: DATA = 8'h00;
            12'b00101_0111110: DATA = 8'h00;
            12'b00101_0111111: DATA = 8'h00;
            12'b00101_1000000: DATA = 8'h00;
            12'b00101_1000001: DATA = 8'h00;
            12'b00101_1000010: DATA = 8'h00;
            12'b00101_1000011: DATA = 8'h00;
            12'b00101_1000100: DATA = 8'h00;
            12'b00101_1000101: DATA = 8'h00;
            12'b00101_1000110: DATA = 8'h00;
            12'b00101_1000111: DATA = 8'h00;
            12'b00101_1001000: DATA = 8'h00;
            12'b00101_1001001: DATA = 8'h00;
            12'b00101_1001010: DATA = 8'h00;
            12'b00101_1001011: DATA = 8'h00;
            12'b00101_1001100: DATA = 8'h00;
            12'b00101_1001101: DATA = 8'h00;
            12'b00101_1001110: DATA = 8'h00;
            12'b00101_1001111: DATA = 8'h00;
            // Row 6
            12'b00110_0000000: DATA = 8'h57;
            12'b00110_0000001: DATA = 8'h41;
            12'b00110_0000010: DATA = 8'h56;
            12'b00110_0000011: DATA = 8'h45;
            12'b00110_0000100: DATA = 8'h46;
            12'b00110_0000101: DATA = 8'h4F;
            12'b00110_0000110: DATA = 8'h52;
            12'b00110_0000111: DATA = 8'h4D;
            12'b00110_0001000: DATA = 8'h00;
            12'b00110_0001001: DATA = 8'h00;
            12'b00110_0001010: DATA = 8'h00;
            12'b00110_0001011: DATA = 8'h00;
            12'b00110_0001100: DATA = 8'h00;
            12'b00110_0001101: DATA = 8'h00;
            12'b00110_0001110: DATA = (WAVE1 == 2'b00) ? 8'h53 : (WAVE1 == 2'b01) ? 8'h53 : (WAVE1 == 2'b10) ? 8'h54 : 8'h53;
            12'b00110_0001111: DATA = (WAVE1 == 2'b00) ? 8'h51 : (WAVE1 == 2'b01) ? 8'h41 : (WAVE1 == 2'b10) ? 8'h52 : 8'h49;
            12'b00110_0010000: DATA = (WAVE1 == 2'b00) ? 8'h55 : (WAVE1 == 2'b01) ? 8'h57 : (WAVE1 == 2'b10) ? 8'h49 : 8'h4E;
            12'b00110_0010001: DATA = (WAVE1 == 2'b00) ? 8'h41 : (WAVE1 == 2'b01) ? 8'h54 : (WAVE1 == 2'b10) ? 8'h41 : 8'h45;
            12'b00110_0010010: DATA = (WAVE1 == 2'b00) ? 8'h52 : (WAVE1 == 2'b01) ? 8'h4F : (WAVE1 == 2'b10) ? 8'h4E : 8'h00;
            12'b00110_0010011: DATA = (WAVE1 == 2'b00) ? 8'h45 : (WAVE1 == 2'b01) ? 8'h4F : (WAVE1 == 2'b10) ? 8'h47 : 8'h00;
            12'b00110_0010100: DATA = (WAVE1 == 2'b00) ? 8'h00 : (WAVE1 == 2'b01) ? 8'h54 : (WAVE1 == 2'b10) ? 8'h4C : 8'h00;
            12'b00110_0010101: DATA = (WAVE1 == 2'b00) ? 8'h00 : (WAVE1 == 2'b01) ? 8'h48 : (WAVE1 == 2'b10) ? 8'h45 : 8'h00;
            12'b00110_0010110: DATA = 8'h00;
            12'b00110_0010111: DATA = 8'h00;
            12'b00110_0011000: DATA = 8'h00;
            12'b00110_0011001: DATA = 8'h00;
            12'b00110_0011010: DATA = 8'h00;
            12'b00110_0011011: DATA = 8'h00;
            12'b00110_0011100: DATA = 8'hC6;
            12'b00110_0011101: DATA = (FORM1 == 2'b10 && WAVE1 == 2'b00) ? 8'hA3 : (FORM1 == 2'b10 && WAVE1 == 2'b01) ? 8'hE7 : (FORM1 == 2'b10 && WAVE1 == 2'b10) ? 8'hB7 : (FORM1 == 2'b10 && WAVE1 == 2'b11) ? 8'h8F : 8'h00;
            12'b00110_0011110: DATA = (FORM1 == 2'b10 && WAVE1 == 2'b00) ? 8'hA4 : (FORM1 == 2'b10 && WAVE1 == 2'b01) ? 8'hE8 : (FORM1 == 2'b10 && WAVE1 == 2'b10) ? 8'hB8 : (FORM1 == 2'b10 && WAVE1 == 2'b11) ? 8'h90 : 8'h00;
            12'b00110_0011111: DATA = (FORM1 == 2'b10 && WAVE1 == 2'b00) ? 8'hA5 : (FORM1 == 2'b10 && WAVE1 == 2'b01) ? 8'hE9 : (FORM1 == 2'b10 && WAVE1 == 2'b10) ? 8'hB9 : (FORM1 == 2'b10 && WAVE1 == 2'b11) ? 8'h91 : 8'h00;
            12'b00110_0100000: DATA = (FORM1 == 2'b10 && WAVE1 == 2'b00) ? 8'hA6 : (FORM1 == 2'b10 && WAVE1 == 2'b01) ? 8'hEA : (FORM1 == 2'b10 && WAVE1 == 2'b10) ? 8'hBA : (FORM1 == 2'b10 && WAVE1 == 2'b11) ? 8'h92 : 8'h00;
            12'b00110_0100001: DATA = (FORM1 == 2'b10 && WAVE1 == 2'b00) ? 8'hA7 : (FORM1 == 2'b10 && WAVE1 == 2'b01) ? 8'hEB : (FORM1 == 2'b10 && WAVE1 == 2'b10) ? 8'hBB : (FORM1 == 2'b10 && WAVE1 == 2'b11) ? 8'h93 : 8'h00;
            12'b00110_0100010: DATA = (FORM1 == 2'b01) ? 8'h00 : (FORM1 == 2'b00 && WAVE1 == 2'b00) ? 8'hA3 : (FORM1 == 2'b00 && WAVE1 == 2'b01) ? 8'hCF : (FORM1 == 2'b00 && WAVE1 == 2'b10) ? 8'hB7 : (FORM1 == 2'b00 && WAVE1 == 2'b11) ? 8'h8F : 8'h00;
            12'b00110_0100011: DATA = (FORM1 == 2'b01) ? 8'h00 : (FORM1 == 2'b00 && WAVE1 == 2'b00) ? 8'hA4 : (FORM1 == 2'b00 && WAVE1 == 2'b01) ? 8'hD0 : (FORM1 == 2'b00 && WAVE1 == 2'b10) ? 8'hB8 : (FORM1 == 2'b00 && WAVE1 == 2'b11) ? 8'h90 : 8'h00;
            12'b00110_0100100: DATA = (FORM1 == 2'b01) ? 8'h00 : (FORM1 == 2'b00 && WAVE1 == 2'b00) ? 8'hA5 : (FORM1 == 2'b00 && WAVE1 == 2'b01) ? 8'hD1 : (FORM1 == 2'b00 && WAVE1 == 2'b10) ? 8'hB9 : (FORM1 == 2'b00 && WAVE1 == 2'b11) ? 8'h91 : 8'h00;
            12'b00110_0100101: DATA = (FORM1 == 2'b01) ? 8'h00 : (FORM1 == 2'b00 && WAVE1 == 2'b00) ? 8'hA6 : (FORM1 == 2'b00 && WAVE1 == 2'b01) ? 8'hD2 : (FORM1 == 2'b00 && WAVE1 == 2'b10) ? 8'hBA : (FORM1 == 2'b00 && WAVE1 == 2'b11) ? 8'h92 : 8'h00;
            12'b00110_0100110: DATA = (FORM1 == 2'b01) ? 8'h00 : (FORM1 == 2'b00 && WAVE1 == 2'b00) ? 8'hA7 : (FORM1 == 2'b00 && WAVE1 == 2'b01) ? 8'hD3 : (FORM1 == 2'b00 && WAVE1 == 2'b10) ? 8'hBB : (FORM1 == 2'b00 && WAVE1 == 2'b11) ? 8'h93 : 8'h00;
            12'b00110_0100111: DATA = 8'hC7;
            12'b00110_0101000: DATA = 8'h00;
            12'b00110_0101001: DATA = 8'h00;
            12'b00110_0101010: DATA = 8'h00;
            12'b00110_0101011: DATA = 8'h00;
            12'b00110_0101100: DATA = 8'h00;
            12'b00110_0101101: DATA = 8'h00;
            12'b00110_0101110: DATA = 8'h00;
            12'b00110_0101111: DATA = 8'h00;
            12'b00110_0110000: DATA = 8'h00;
            12'b00110_0110001: DATA = 8'h00;
            12'b00110_0110010: DATA = 8'h00;
            12'b00110_0110011: DATA = 8'h00;
            12'b00110_0110100: DATA = 8'h00;
            12'b00110_0110101: DATA = 8'h00;
            12'b00110_0110110: DATA = 8'h00;
            12'b00110_0110111: DATA = 8'h00;
            12'b00110_0111000: DATA = 8'h00;
            12'b00110_0111001: DATA = 8'h00;
            12'b00110_0111010: DATA = 8'h00;
            12'b00110_0111011: DATA = 8'h00;
            12'b00110_0111100: DATA = 8'h00;
            12'b00110_0111101: DATA = 8'h00;
            12'b00110_0111110: DATA = 8'h00;
            12'b00110_0111111: DATA = 8'h00;
            12'b00110_1000000: DATA = 8'h00;
            12'b00110_1000001: DATA = 8'h00;
            12'b00110_1000010: DATA = 8'h00;
            12'b00110_1000011: DATA = 8'h00;
            12'b00110_1000100: DATA = 8'h00;
            12'b00110_1000101: DATA = 8'h00;
            12'b00110_1000110: DATA = 8'h00;
            12'b00110_1000111: DATA = 8'h00;
            12'b00110_1001000: DATA = 8'h00;
            12'b00110_1001001: DATA = 8'h00;
            12'b00110_1001010: DATA = 8'h00;
            12'b00110_1001011: DATA = 8'h00;
            12'b00110_1001100: DATA = 8'h00;
            12'b00110_1001101: DATA = 8'h00;
            12'b00110_1001110: DATA = 8'h00;
            12'b00110_1001111: DATA = 8'h00;
            // Row 7
            12'b00111_0000000: DATA = 8'h4D;
            12'b00111_0000001: DATA = 8'h4F;
            12'b00111_0000010: DATA = 8'h44;
            12'b00111_0000011: DATA = 8'h45;
            12'b00111_0000100: DATA = 8'h00;
            12'b00111_0000101: DATA = 8'h00;
            12'b00111_0000110: DATA = 8'h00;
            12'b00111_0000111: DATA = 8'h00;
            12'b00111_0001000: DATA = 8'h00;
            12'b00111_0001001: DATA = 8'h00;
            12'b00111_0001010: DATA = 8'h00;
            12'b00111_0001011: DATA = 8'h00;
            12'b00111_0001100: DATA = 8'h00;
            12'b00111_0001101: DATA = 8'h00;
            12'b00111_0001110: DATA = (FORM1 == 2'b00) ? 8'h4E : (FORM1 == 2'b01) ? 8'h48 : (FORM1 == 2'b10) ? 8'h52 : 8'h46;
            12'b00111_0001111: DATA = (FORM1 == 2'b00) ? 8'h4F : (FORM1 == 2'b01) ? 8'h41 : (FORM1 == 2'b10) ? 8'h45 : 8'h55;
            12'b00111_0010000: DATA = (FORM1 == 2'b00) ? 8'h52 : (FORM1 == 2'b01) ? 8'h4C : (FORM1 == 2'b10) ? 8'h56 : 8'h4C;
            12'b00111_0010001: DATA = (FORM1 == 2'b00) ? 8'h4D : (FORM1 == 2'b01) ? 8'h46 : (FORM1 == 2'b10) ? 8'h45 : 8'h4C;
            12'b00111_0010010: DATA = (FORM1 == 2'b00) ? 8'h41 : (FORM1 == 2'b01) ? 8'h2D : (FORM1 == 2'b10) ? 8'h52 : 8'h2D;
            12'b00111_0010011: DATA = (FORM1 == 2'b00) ? 8'h4C : (FORM1 == 2'b01) ? 8'h57 : (FORM1 == 2'b10) ? 8'h53 : 8'h57;
            12'b00111_0010100: DATA = (FORM1 == 2'b00) ? 8'h00 : (FORM1 == 2'b01) ? 8'h41 : (FORM1 == 2'b10) ? 8'h45 : 8'h41;
            12'b00111_0010101: DATA = (FORM1 == 2'b00) ? 8'h00 : (FORM1 == 2'b01) ? 8'h56 : (FORM1 == 2'b10) ? 8'h44 : 8'h56;
            12'b00111_0010110: DATA = (FORM1 == 2'b00) ? 8'h00 : (FORM1 == 2'b01) ? 8'h45 : (FORM1 == 2'b10) ? 8'h00 : 8'h45;
            12'b00111_0010111: DATA = 8'h00;
            12'b00111_0011000: DATA = 8'h00;
            12'b00111_0011001: DATA = 8'h00;
            12'b00111_0011010: DATA = 8'h00;
            12'b00111_0011011: DATA = 8'h00;
            12'b00111_0011100: DATA = 8'hD6;
            12'b00111_0011101: DATA = 8'hC9;
            12'b00111_0011110: DATA = 8'hC9;
            12'b00111_0011111: DATA = 8'hC9;
            12'b00111_0100000: DATA = 8'hC9;
            12'b00111_0100001: DATA = 8'hC9;
            12'b00111_0100010: DATA = 8'hC9;
            12'b00111_0100011: DATA = 8'hC9;
            12'b00111_0100100: DATA = 8'hC9;
            12'b00111_0100101: DATA = 8'hC9;
            12'b00111_0100110: DATA = 8'hC9;
            12'b00111_0100111: DATA = 8'hD7;
            12'b00111_0101000: DATA = 8'h00;
            12'b00111_0101001: DATA = 8'h00;
            12'b00111_0101010: DATA = 8'h00;
            12'b00111_0101011: DATA = 8'h00;
            12'b00111_0101100: DATA = 8'h00;
            12'b00111_0101101: DATA = 8'h00;
            12'b00111_0101110: DATA = 8'h00;
            12'b00111_0101111: DATA = 8'h00;
            12'b00111_0110000: DATA = 8'h00;
            12'b00111_0110001: DATA = 8'h00;
            12'b00111_0110010: DATA = 8'h00;
            12'b00111_0110011: DATA = 8'h00;
            12'b00111_0110100: DATA = 8'h00;
            12'b00111_0110101: DATA = 8'h00;
            12'b00111_0110110: DATA = 8'h00;
            12'b00111_0110111: DATA = 8'h00;
            12'b00111_0111000: DATA = 8'h00;
            12'b00111_0111001: DATA = 8'h00;
            12'b00111_0111010: DATA = 8'h00;
            12'b00111_0111011: DATA = 8'h00;
            12'b00111_0111100: DATA = 8'h00;
            12'b00111_0111101: DATA = 8'h00;
            12'b00111_0111110: DATA = 8'h00;
            12'b00111_0111111: DATA = 8'h00;
            12'b00111_1000000: DATA = 8'h00;
            12'b00111_1000001: DATA = 8'h00;
            12'b00111_1000010: DATA = 8'h00;
            12'b00111_1000011: DATA = 8'h00;
            12'b00111_1000100: DATA = 8'h00;
            12'b00111_1000101: DATA = 8'h00;
            12'b00111_1000110: DATA = 8'h00;
            12'b00111_1000111: DATA = 8'h00;
            12'b00111_1001000: DATA = 8'h00;
            12'b00111_1001001: DATA = 8'h00;
            12'b00111_1001010: DATA = 8'h00;
            12'b00111_1001011: DATA = 8'h00;
            12'b00111_1001100: DATA = 8'h00;
            12'b00111_1001101: DATA = 8'h00;
            12'b00111_1001110: DATA = 8'h00;
            12'b00111_1001111: DATA = 8'h00;
            // Row 8
            12'b01000_0000000: DATA = 8'h00;
            12'b01000_0000001: DATA = 8'h00;
            12'b01000_0000010: DATA = 8'h00;
            12'b01000_0000011: DATA = 8'h00;
            12'b01000_0000100: DATA = 8'h00;
            12'b01000_0000101: DATA = 8'h00;
            12'b01000_0000110: DATA = 8'h00;
            12'b01000_0000111: DATA = 8'h00;
            12'b01000_0001000: DATA = 8'h00;
            12'b01000_0001001: DATA = 8'h00;
            12'b01000_0001010: DATA = 8'h00;
            12'b01000_0001011: DATA = 8'h00;
            12'b01000_0001100: DATA = 8'h00;
            12'b01000_0001101: DATA = 8'h00;
            12'b01000_0001110: DATA = 8'h00;
            12'b01000_0001111: DATA = 8'h00;
            12'b01000_0010000: DATA = 8'h00;
            12'b01000_0010001: DATA = 8'h00;
            12'b01000_0010010: DATA = 8'h00;
            12'b01000_0010011: DATA = 8'h00;
            12'b01000_0010100: DATA = 8'h00;
            12'b01000_0010101: DATA = 8'h00;
            12'b01000_0010110: DATA = 8'h00;
            12'b01000_0010111: DATA = 8'h00;
            12'b01000_0011000: DATA = 8'h00;
            12'b01000_0011001: DATA = 8'h00;
            12'b01000_0011010: DATA = 8'h00;
            12'b01000_0011011: DATA = 8'h00;
            12'b01000_0011100: DATA = 8'h00;
            12'b01000_0011101: DATA = 8'h00;
            12'b01000_0011110: DATA = 8'h00;
            12'b01000_0011111: DATA = 8'h00;
            12'b01000_0100000: DATA = 8'h00;
            12'b01000_0100001: DATA = 8'h00;
            12'b01000_0100010: DATA = 8'h00;
            12'b01000_0100011: DATA = 8'h00;
            12'b01000_0100100: DATA = 8'h00;
            12'b01000_0100101: DATA = 8'h00;
            12'b01000_0100110: DATA = 8'h00;
            12'b01000_0100111: DATA = 8'h00;
            12'b01000_0101000: DATA = 8'h00;
            12'b01000_0101001: DATA = 8'h00;
            12'b01000_0101010: DATA = 8'h00;
            12'b01000_0101011: DATA = 8'h00;
            12'b01000_0101100: DATA = 8'h00;
            12'b01000_0101101: DATA = 8'h00;
            12'b01000_0101110: DATA = 8'h00;
            12'b01000_0101111: DATA = 8'h00;
            12'b01000_0110000: DATA = 8'h00;
            12'b01000_0110001: DATA = 8'h00;
            12'b01000_0110010: DATA = 8'h00;
            12'b01000_0110011: DATA = 8'h00;
            12'b01000_0110100: DATA = 8'h00;
            12'b01000_0110101: DATA = 8'h00;
            12'b01000_0110110: DATA = 8'h00;
            12'b01000_0110111: DATA = 8'h00;
            12'b01000_0111000: DATA = 8'h00;
            12'b01000_0111001: DATA = 8'h00;
            12'b01000_0111010: DATA = 8'h00;
            12'b01000_0111011: DATA = 8'h00;
            12'b01000_0111100: DATA = 8'h00;
            12'b01000_0111101: DATA = 8'h00;
            12'b01000_0111110: DATA = 8'h00;
            12'b01000_0111111: DATA = 8'h00;
            12'b01000_1000000: DATA = 8'h00;
            12'b01000_1000001: DATA = 8'h00;
            12'b01000_1000010: DATA = 8'h00;
            12'b01000_1000011: DATA = 8'h00;
            12'b01000_1000100: DATA = 8'h00;
            12'b01000_1000101: DATA = 8'h00;
            12'b01000_1000110: DATA = 8'h00;
            12'b01000_1000111: DATA = 8'h00;
            12'b01000_1001000: DATA = 8'h00;
            12'b01000_1001001: DATA = 8'h00;
            12'b01000_1001010: DATA = 8'h00;
            12'b01000_1001011: DATA = 8'h00;
            12'b01000_1001100: DATA = 8'h00;
            12'b01000_1001101: DATA = 8'h00;
            12'b01000_1001110: DATA = 8'h00;
            12'b01000_1001111: DATA = 8'h00;
            // Row 9
            12'b01001_0000000: DATA = 8'h43;
            12'b01001_0000001: DATA = 8'h48;
            12'b01001_0000010: DATA = 8'h41;
            12'b01001_0000011: DATA = 8'h4E;
            12'b01001_0000100: DATA = 8'h4E;
            12'b01001_0000101: DATA = 8'h45;
            12'b01001_0000110: DATA = 8'h4C;
            12'b01001_0000111: DATA = 8'h00;
            12'b01001_0001000: DATA = 8'h32;
            12'b01001_0001001: DATA = 8'h00;
            12'b01001_0001010: DATA = (CHANNEL == 1) ? 8'h3C : 8'h00;
            12'b01001_0001011: DATA = 8'h00;
            12'b01001_0001100: DATA = (CHANNEL == 1 && DC == 1) ? 8'h44 : 8'h00;
            12'b01001_0001101: DATA = (CHANNEL == 1 && DC == 1) ? 8'h43 : 8'h00;
            12'b01001_0001110: DATA = 8'h00;
            12'b01001_0001111: DATA = 8'h00;
            12'b01001_0010000: DATA = 8'h00;
            12'b01001_0010001: DATA = 8'h00;
            12'b01001_0010010: DATA = 8'h00;
            12'b01001_0010011: DATA = 8'h00;
            12'b01001_0010100: DATA = 8'h00;
            12'b01001_0010101: DATA = 8'h00;
            12'b01001_0010110: DATA = 8'h00;
            12'b01001_0010111: DATA = 8'h00;
            12'b01001_0011000: DATA = 8'h00;
            12'b01001_0011001: DATA = 8'h00;
            12'b01001_0011010: DATA = 8'h00;
            12'b01001_0011011: DATA = 8'h00;
            12'b01001_0011100: DATA = 8'hD4;
            12'b01001_0011101: DATA = 8'hC8;
            12'b01001_0011110: DATA = 8'hC8;
            12'b01001_0011111: DATA = 8'hC8;
            12'b01001_0100000: DATA = 8'hC8;
            12'b01001_0100001: DATA = 8'hC8;
            12'b01001_0100010: DATA = 8'hC8;
            12'b01001_0100011: DATA = 8'hC8;
            12'b01001_0100100: DATA = 8'hC8;
            12'b01001_0100101: DATA = 8'hC8;
            12'b01001_0100110: DATA = 8'hC8;
            12'b01001_0100111: DATA = 8'hD5;
            12'b01001_0101000: DATA = 8'h00;
            12'b01001_0101001: DATA = 8'h00;
            12'b01001_0101010: DATA = 8'h00;
            12'b01001_0101011: DATA = 8'h00;
            12'b01001_0101100: DATA = 8'h00;
            12'b01001_0101101: DATA = 8'h00;
            12'b01001_0101110: DATA = 8'h00;
            12'b01001_0101111: DATA = 8'h00;
            12'b01001_0110000: DATA = 8'h00;
            12'b01001_0110001: DATA = 8'h00;
            12'b01001_0110010: DATA = 8'h00;
            12'b01001_0110011: DATA = 8'h00;
            12'b01001_0110100: DATA = 8'h00;
            12'b01001_0110101: DATA = 8'h00;
            12'b01001_0110110: DATA = 8'h00;
            12'b01001_0110111: DATA = 8'h00;
            12'b01001_0111000: DATA = 8'h00;
            12'b01001_0111001: DATA = 8'h00;
            12'b01001_0111010: DATA = 8'h00;
            12'b01001_0111011: DATA = 8'h00;
            12'b01001_0111100: DATA = 8'h00;
            12'b01001_0111101: DATA = 8'h00;
            12'b01001_0111110: DATA = 8'h00;
            12'b01001_0111111: DATA = 8'h00;
            12'b01001_1000000: DATA = 8'h00;
            12'b01001_1000001: DATA = 8'h00;
            12'b01001_1000010: DATA = 8'h00;
            12'b01001_1000011: DATA = 8'h00;
            12'b01001_1000100: DATA = 8'h00;
            12'b01001_1000101: DATA = 8'h00;
            12'b01001_1000110: DATA = 8'h00;
            12'b01001_1000111: DATA = 8'h00;
            12'b01001_1001000: DATA = 8'h00;
            12'b01001_1001001: DATA = 8'h00;
            12'b01001_1001010: DATA = 8'h00;
            12'b01001_1001011: DATA = 8'h00;
            12'b01001_1001100: DATA = 8'h00;
            12'b01001_1001101: DATA = 8'h00;
            12'b01001_1001110: DATA = 8'h00;
            12'b01001_1001111: DATA = 8'h00;
            // Row 10
            12'b01010_0000000: DATA = 8'h46;
            12'b01010_0000001: DATA = 8'h52;
            12'b01010_0000010: DATA = 8'h45;
            12'b01010_0000011: DATA = 8'h51;
            12'b01010_0000100: DATA = 8'h55;
            12'b01010_0000101: DATA = 8'h45;
            12'b01010_0000110: DATA = 8'h4E;
            12'b01010_0000111: DATA = 8'h43;
            12'b01010_0001000: DATA = 8'h59;
            12'b01010_0001001: DATA = 8'h00;
            12'b01010_0001010: DATA = 8'h00;
            12'b01010_0001011: DATA = 8'h00;
            12'b01010_0001100: DATA = 8'h00;
            12'b01010_0001101: DATA = 8'h00;
            12'b01010_0001110: DATA = FREQ2[39:32];
            12'b01010_0001111: DATA = FREQ2[31:24];
            12'b01010_0010000: DATA = FREQ2[23:16];
            12'b01010_0010001: DATA = FREQ2[15:8];
            12'b01010_0010010: DATA = FREQ2[7:0];
            12'b01010_0010011: DATA = 8'h00;
            12'b01010_0010100: DATA = 8'h00;
            12'b01010_0010101: DATA = 8'h00;
            12'b01010_0010110: DATA = 8'h00;
            12'b01010_0010111: DATA = 8'h00;
            12'b01010_0011000: DATA = 8'h00;
            12'b01010_0011001: DATA = 8'h00;
            12'b01010_0011010: DATA = 8'h00;
            12'b01010_0011011: DATA = 8'h00;
            12'b01010_0011100: DATA = 8'hC6;
            12'b01010_0011101: DATA = (FORM2 == 2'b10) ? 8'h00 : (WAVE2 == 2'b00) ? 8'h94 : (WAVE2 == 2'b01) ? 8'hBC : (WAVE2 == 2'b10) ? 8'hA8 : 8'h80;
            12'b01010_0011110: DATA = (FORM2 == 2'b10) ? 8'h00 : (WAVE2 == 2'b00) ? 8'h95 : (WAVE2 == 2'b01) ? 8'hBD : (WAVE2 == 2'b10) ? 8'hA9 : 8'h81;
            12'b01010_0011111: DATA = (FORM2 == 2'b10) ? 8'h00 : (WAVE2 == 2'b00) ? 8'h96 : (WAVE2 == 2'b01) ? 8'hBE : (WAVE2 == 2'b10) ? 8'hAA : 8'h82;
            12'b01010_0100000: DATA = (FORM2 == 2'b10) ? 8'h00 : (WAVE2 == 2'b00) ? 8'h97 : (WAVE2 == 2'b01) ? 8'hBF : (WAVE2 == 2'b10) ? 8'hAB : 8'h83;
            12'b01010_0100001: DATA = (FORM2 == 2'b10) ? 8'h00 : (WAVE2 == 2'b00) ? 8'h98 : (WAVE2 == 2'b01) ? 8'hC0 : (WAVE2 == 2'b10) ? 8'hAC : 8'h84;
            12'b01010_0100010: DATA = (FORM2 == 2'b00) ? 8'h00 : (FORM2 == 2'b01) ? 8'h00 : (WAVE2 == 2'b00) ? 8'h94 : (WAVE2 == 2'b01) ? 8'hD8 : (WAVE2 == 2'b10) ? 8'hA8 : 8'h80;
            12'b01010_0100011: DATA = (FORM2 == 2'b00) ? 8'h00 : (FORM2 == 2'b01) ? 8'h00 : (WAVE2 == 2'b00) ? 8'h95 : (WAVE2 == 2'b01) ? 8'hD9 : (WAVE2 == 2'b10) ? 8'hA9 : 8'h81;
            12'b01010_0100100: DATA = (FORM2 == 2'b00) ? 8'h00 : (FORM2 == 2'b01) ? 8'h00 : (WAVE2 == 2'b00) ? 8'h96 : (WAVE2 == 2'b01) ? 8'hDA : (WAVE2 == 2'b10) ? 8'hAA : 8'h82;
            12'b01010_0100101: DATA = (FORM2 == 2'b00) ? 8'h00 : (FORM2 == 2'b01) ? 8'h00 : (WAVE2 == 2'b00) ? 8'h97 : (WAVE2 == 2'b01) ? 8'hDB : (WAVE2 == 2'b10) ? 8'hAB : 8'h83;
            12'b01010_0100110: DATA = (FORM2 == 2'b00) ? 8'h00 : (FORM2 == 2'b01) ? 8'h00 : (WAVE2 == 2'b00) ? 8'h98 : (WAVE2 == 2'b01) ? 8'hDC : (WAVE2 == 2'b10) ? 8'hAC : 8'h84;
            12'b01010_0100111: DATA = 8'hC7;
            12'b01010_0101000: DATA = 8'h00;
            12'b01010_0101001: DATA = 8'h00;
            12'b01010_0101010: DATA = 8'h00;
            12'b01010_0101011: DATA = 8'h00;
            12'b01010_0101100: DATA = 8'h00;
            12'b01010_0101101: DATA = 8'h00;
            12'b01010_0101110: DATA = 8'h00;
            12'b01010_0101111: DATA = 8'h00;
            12'b01010_0110000: DATA = 8'h00;
            12'b01010_0110001: DATA = 8'h00;
            12'b01010_0110010: DATA = 8'h00;
            12'b01010_0110011: DATA = 8'h00;
            12'b01010_0110100: DATA = 8'h00;
            12'b01010_0110101: DATA = 8'h00;
            12'b01010_0110110: DATA = 8'h00;
            12'b01010_0110111: DATA = 8'h00;
            12'b01010_0111000: DATA = 8'h00;
            12'b01010_0111001: DATA = 8'h00;
            12'b01010_0111010: DATA = 8'h00;
            12'b01010_0111011: DATA = 8'h00;
            12'b01010_0111100: DATA = 8'h00;
            12'b01010_0111101: DATA = 8'h00;
            12'b01010_0111110: DATA = 8'h00;
            12'b01010_0111111: DATA = 8'h00;
            12'b01010_1000000: DATA = 8'h00;
            12'b01010_1000001: DATA = 8'h00;
            12'b01010_1000010: DATA = 8'h00;
            12'b01010_1000011: DATA = 8'h00;
            12'b01010_1000100: DATA = 8'h00;
            12'b01010_1000101: DATA = 8'h00;
            12'b01010_1000110: DATA = 8'h00;
            12'b01010_1000111: DATA = 8'h00;
            12'b01010_1001000: DATA = 8'h00;
            12'b01010_1001001: DATA = 8'h00;
            12'b01010_1001010: DATA = 8'h00;
            12'b01010_1001011: DATA = 8'h00;
            12'b01010_1001100: DATA = 8'h00;
            12'b01010_1001101: DATA = 8'h00;
            12'b01010_1001110: DATA = 8'h00;
            12'b01010_1001111: DATA = 8'h00;
            // Row 11
            12'b01011_0000000: DATA = 8'h4D;
            12'b01011_0000001: DATA = 8'h41;
            12'b01011_0000010: DATA = 8'h58;
            12'b01011_0000011: DATA = 8'h00;
            12'b01011_0000100: DATA = 8'h41;
            12'b01011_0000101: DATA = 8'h4D;
            12'b01011_0000110: DATA = 8'h50;
            12'b01011_0000111: DATA = 8'h4C;
            12'b01011_0001000: DATA = 8'h49;
            12'b01011_0001001: DATA = 8'h54;
            12'b01011_0001010: DATA = 8'h55;
            12'b01011_0001011: DATA = 8'h44;
            12'b01011_0001100: DATA = 8'h45;
            12'b01011_0001101: DATA = 8'h00;
            12'b01011_0001110: DATA = MAX_AMP2[31:24];
            12'b01011_0001111: DATA = (AMP_MODE == 1) ? MAX_AMP2[23:16] : 8'h2E;
            12'b01011_0010000: DATA = (AMP_MODE == 1) ? MAX_AMP2[15:8] : MAX_AMP2[23:16];
            12'b01011_0010001: DATA = (AMP_MODE == 1) ? MAX_AMP2[7:0] : MAX_AMP2[15:8];
            12'b01011_0010010: DATA = (AMP_MODE == 1) ? 8'h00 : MAX_AMP2[7:0];
            12'b01011_0010011: DATA = 8'h00;
            12'b01011_0010100: DATA = 8'h00;
            12'b01011_0010101: DATA = 8'h00;
            12'b01011_0010110: DATA = 8'h00;
            12'b01011_0010111: DATA = 8'h00;
            12'b01011_0011000: DATA = 8'h00;
            12'b01011_0011001: DATA = 8'h00;
            12'b01011_0011010: DATA = 8'h00;
            12'b01011_0011011: DATA = 8'h00;
            12'b01011_0011100: DATA = 8'hC6;
            12'b01011_0011101: DATA = (FORM2 == 2'b10) ? 8'h00 : (WAVE2 == 2'b00) ? 8'h99 : (WAVE2 == 2'b01) ? 8'hC1 : (WAVE2 == 2'b10) ? 8'hAD : 8'h85;
            12'b01011_0011110: DATA = (FORM2 == 2'b10) ? 8'h00 : (WAVE2 == 2'b00) ? 8'h9A : (WAVE2 == 2'b01) ? 8'hC2 : (WAVE2 == 2'b10) ? 8'hAE : 8'h86;
            12'b01011_0011111: DATA = (FORM2 == 2'b10) ? 8'h00 : (WAVE2 == 2'b00) ? 8'h9B : (WAVE2 == 2'b01) ? 8'hC3 : (WAVE2 == 2'b10) ? 8'hAF : 8'h87;
            12'b01011_0100000: DATA = (FORM2 == 2'b10) ? 8'h00 : (WAVE2 == 2'b00) ? 8'h9C : (WAVE2 == 2'b01) ? 8'hC4 : (WAVE2 == 2'b10) ? 8'hB0 : 8'h88;
            12'b01011_0100001: DATA = (FORM2 == 2'b10) ? 8'h00 : (WAVE2 == 2'b00) ? 8'h9D : (WAVE2 == 2'b01) ? 8'hC5 : (WAVE2 == 2'b10) ? 8'hB1 : 8'h89;
            12'b01011_0100010: DATA = (FORM2 == 2'b00) ? 8'h00 : (FORM2 == 2'b01) ? 8'h00 : (WAVE2 == 2'b00) ? 8'h99 : (WAVE2 == 2'b01) ? 8'hDD: (WAVE2 == 2'b10) ? 8'hAD : 8'h85;
            12'b01011_0100011: DATA = (FORM2 == 2'b00) ? 8'h00 : (FORM2 == 2'b01) ? 8'h00 : (WAVE2 == 2'b00) ? 8'h9A : (WAVE2 == 2'b01) ? 8'hDE : (WAVE2 == 2'b10) ? 8'hAE : 8'h86;
            12'b01011_0100100: DATA = (FORM2 == 2'b00) ? 8'h00 : (FORM2 == 2'b01) ? 8'h00 : (WAVE2 == 2'b00) ? 8'h9B : (WAVE2 == 2'b01) ? 8'hDF : (WAVE2 == 2'b10) ? 8'hAF : 8'h87;
            12'b01011_0100101: DATA = (FORM2 == 2'b00) ? 8'h00 : (FORM2 == 2'b01) ? 8'h00 : (WAVE2 == 2'b00) ? 8'h9C : (WAVE2 == 2'b01) ? 8'hE0 : (WAVE2 == 2'b10) ? 8'hB0 : 8'h88;
            12'b01011_0100110: DATA = (FORM2 == 2'b00) ? 8'h00 : (FORM2 == 2'b01) ? 8'h00 : (WAVE2 == 2'b00) ? 8'h9D : (WAVE2 == 2'b01) ? 8'hE1 : (WAVE2 == 2'b10) ? 8'hB1 : 8'h89;
            12'b01011_0100111: DATA = 8'hC7;
            12'b01011_0101000: DATA = 8'h00;
            12'b01011_0101001: DATA = 8'h00;
            12'b01011_0101010: DATA = 8'h00;
            12'b01011_0101011: DATA = 8'h00;
            12'b01011_0101100: DATA = 8'h00;
            12'b01011_0101101: DATA = 8'h00;
            12'b01011_0101110: DATA = 8'h00;
            12'b01011_0101111: DATA = 8'h00;
            12'b01011_0110000: DATA = 8'h00;
            12'b01011_0110001: DATA = 8'h00;
            12'b01011_0110010: DATA = 8'h00;
            12'b01011_0110011: DATA = 8'h00;
            12'b01011_0110100: DATA = 8'h00;
            12'b01011_0110101: DATA = 8'h00;
            12'b01011_0110110: DATA = 8'h00;
            12'b01011_0110111: DATA = 8'h00;
            12'b01011_0111000: DATA = 8'h00;
            12'b01011_0111001: DATA = 8'h00;
            12'b01011_0111010: DATA = 8'h00;
            12'b01011_0111011: DATA = 8'h00;
            12'b01011_0111100: DATA = 8'h00;
            12'b01011_0111101: DATA = 8'h00;
            12'b01011_0111110: DATA = 8'h00;
            12'b01011_0111111: DATA = 8'h00;
            12'b01011_1000000: DATA = 8'h00;
            12'b01011_1000001: DATA = 8'h00;
            12'b01011_1000010: DATA = 8'h00;
            12'b01011_1000011: DATA = 8'h00;
            12'b01011_1000100: DATA = 8'h00;
            12'b01011_1000101: DATA = 8'h00;
            12'b01011_1000110: DATA = 8'h00;
            12'b01011_1000111: DATA = 8'h00;
            12'b01011_1001000: DATA = 8'h00;
            12'b01011_1001001: DATA = 8'h00;
            12'b01011_1001010: DATA = 8'h00;
            12'b01011_1001011: DATA = 8'h00;
            12'b01011_1001100: DATA = 8'h00;
            12'b01011_1001101: DATA = 8'h00;
            12'b01011_1001110: DATA = 8'h00;
            12'b01011_1001111: DATA = 8'h00;
            // Row 12
            12'b01100_0000000: DATA = 8'h4D;
            12'b01100_0000001: DATA = 8'h49;
            12'b01100_0000010: DATA = 8'h4E;
            12'b01100_0000011: DATA = 8'h00;
            12'b01100_0000100: DATA = 8'h41;
            12'b01100_0000101: DATA = 8'h4D;
            12'b01100_0000110: DATA = 8'h50;
            12'b01100_0000111: DATA = 8'h4C;
            12'b01100_0001000: DATA = 8'h49;
            12'b01100_0001001: DATA = 8'h54;
            12'b01100_0001010: DATA = 8'h55;
            12'b01100_0001011: DATA = 8'h44;
            12'b01100_0001100: DATA = 8'h45;
            12'b01100_0001101: DATA = 8'h00;
            12'b01100_0001110: DATA = MIN_AMP2[31:24];
            12'b01100_0001111: DATA = (AMP_MODE == 1) ? MIN_AMP2[23:16] : 8'h2E;
            12'b01100_0010000: DATA = (AMP_MODE == 1) ? MIN_AMP2[15:8] : MIN_AMP2[23:16];
            12'b01100_0010001: DATA = (AMP_MODE == 1) ? MIN_AMP2[7:0] : MIN_AMP2[15:8];
            12'b01100_0010010: DATA = (AMP_MODE == 1) ? 8'h00 : MIN_AMP2[7:0];
            12'b01100_0010011: DATA = 8'h00;
            12'b01100_0010100: DATA = 8'h00;
            12'b01100_0010101: DATA = 8'h00;
            12'b01100_0010110: DATA = 8'h00;
            12'b01100_0010111: DATA = 8'h00;
            12'b01100_0011000: DATA = 8'h00;
            12'b01100_0011001: DATA = 8'h00;
            12'b01100_0011010: DATA = 8'h00;
            12'b01100_0011011: DATA = 8'h00;
            12'b01100_0011100: DATA = 8'hC6;
            12'b01100_0011101: DATA = (FORM2 == 2'b10 && WAVE2 == 2'b00) ? 8'h9E : (FORM2 == 2'b10 && WAVE2 == 2'b01) ? 8'hE2 : (FORM2 == 2'b10 && WAVE2 == 2'b10) ? 8'hB2 : (FORM2 == 2'b10 && WAVE2 == 2'b11) ? 8'h8A : 8'h00;
            12'b01100_0011110: DATA = (FORM2 == 2'b10 && WAVE2 == 2'b00) ? 8'h9F : (FORM2 == 2'b10 && WAVE2 == 2'b01) ? 8'hE3 : (FORM2 == 2'b10 && WAVE2 == 2'b10) ? 8'hB3 : (FORM2 == 2'b10 && WAVE2 == 2'b11) ? 8'h8B : 8'h00;
            12'b01100_0011111: DATA = (FORM2 == 2'b10 && WAVE2 == 2'b00) ? 8'hA0 : (FORM2 == 2'b10 && WAVE2 == 2'b01) ? 8'hE4 : (FORM2 == 2'b10 && WAVE2 == 2'b10) ? 8'hB4 : (FORM2 == 2'b10 && WAVE2 == 2'b11) ? 8'h8C : 8'h00;
            12'b01100_0100000: DATA = (FORM2 == 2'b10 && WAVE2 == 2'b00) ? 8'hA1 : (FORM2 == 2'b10 && WAVE2 == 2'b01) ? 8'hE5 : (FORM2 == 2'b10 && WAVE2 == 2'b10) ? 8'hB5 : (FORM2 == 2'b10 && WAVE2 == 2'b11) ? 8'h8D : 8'h00;
            12'b01100_0100001: DATA = (FORM2 == 2'b10 && WAVE2 == 2'b00) ? 8'hA2 : (FORM2 == 2'b10 && WAVE2 == 2'b01) ? 8'hE6 : (FORM2 == 2'b10 && WAVE2 == 2'b10) ? 8'hB6 : (FORM2 == 2'b10 && WAVE2 == 2'b11) ? 8'h8E : 8'h00;
            12'b01100_0100010: DATA = (FORM2 == 2'b01) ? 8'hC8 : (FORM2 == 2'b00 && WAVE2 == 2'b00) ? 8'h9E : (FORM2 == 2'b00 && WAVE2 == 2'b01) ? 8'hCA : (FORM2 == 2'b00 && WAVE2 == 2'b10) ? 8'hB2 : (FORM2 == 2'b00 && WAVE2 == 2'b11) ? 8'h8A : 8'h00;
            12'b01100_0100011: DATA = (FORM2 == 2'b01) ? 8'hC8 : (FORM2 == 2'b00 && WAVE2 == 2'b00) ? 8'h9F : (FORM2 == 2'b00 && WAVE2 == 2'b01) ? 8'hCB : (FORM2 == 2'b00 && WAVE2 == 2'b10) ? 8'hB3 : (FORM2 == 2'b00 && WAVE2 == 2'b11) ? 8'h8B : 8'h00;
            12'b01100_0100100: DATA = (FORM2 == 2'b01) ? 8'hC8 : (FORM2 == 2'b00 && WAVE2 == 2'b00) ? 8'hA0 : (FORM2 == 2'b00 && WAVE2 == 2'b01) ? 8'hCC : (FORM2 == 2'b00 && WAVE2 == 2'b10) ? 8'hB4 : (FORM2 == 2'b00 && WAVE2 == 2'b11) ? 8'h8C : 8'h00;
            12'b01100_0100101: DATA = (FORM2 == 2'b01) ? 8'hC8 : (FORM2 == 2'b00 && WAVE2 == 2'b00) ? 8'hA1 : (FORM2 == 2'b00 && WAVE2 == 2'b01) ? 8'hCD : (FORM2 == 2'b00 && WAVE2 == 2'b10) ? 8'hB5 : (FORM2 == 2'b00 && WAVE2 == 2'b11) ? 8'h8D : 8'h00;
            12'b01100_0100110: DATA = (FORM2 == 2'b01) ? 8'hC8 : (FORM2 == 2'b00 && WAVE2 == 2'b00) ? 8'hA2 : (FORM2 == 2'b00 && WAVE2 == 2'b01) ? 8'hCE : (FORM2 == 2'b00 && WAVE2 == 2'b10) ? 8'hB6 : (FORM2 == 2'b00 && WAVE2 == 2'b11) ? 8'h8E : 8'h00;
            12'b01100_0100111: DATA = 8'hC7;
            12'b01100_0101000: DATA = 8'h00;
            12'b01100_0101001: DATA = 8'h00;
            12'b01100_0101010: DATA = 8'h00;
            12'b01100_0101011: DATA = 8'h00;
            12'b01100_0101100: DATA = 8'h00;
            12'b01100_0101101: DATA = 8'h00;
            12'b01100_0101110: DATA = 8'h00;
            12'b01100_0101111: DATA = 8'h00;
            12'b01100_0110000: DATA = 8'h00;
            12'b01100_0110001: DATA = 8'h00;
            12'b01100_0110010: DATA = 8'h00;
            12'b01100_0110011: DATA = 8'h00;
            12'b01100_0110100: DATA = 8'h00;
            12'b01100_0110101: DATA = 8'h00;
            12'b01100_0110110: DATA = 8'h00;
            12'b01100_0110111: DATA = 8'h00;
            12'b01100_0111000: DATA = 8'h00;
            12'b01100_0111001: DATA = 8'h00;
            12'b01100_0111010: DATA = 8'h00;
            12'b01100_0111011: DATA = 8'h00;
            12'b01100_0111100: DATA = 8'h00;
            12'b01100_0111101: DATA = 8'h00;
            12'b01100_0111110: DATA = 8'h00;
            12'b01100_0111111: DATA = 8'h00;
            12'b01100_1000000: DATA = 8'h00;
            12'b01100_1000001: DATA = 8'h00;
            12'b01100_1000010: DATA = 8'h00;
            12'b01100_1000011: DATA = 8'h00;
            12'b01100_1000100: DATA = 8'h00;
            12'b01100_1000101: DATA = 8'h00;
            12'b01100_1000110: DATA = 8'h00;
            12'b01100_1000111: DATA = 8'h00;
            12'b01100_1001000: DATA = 8'h00;
            12'b01100_1001001: DATA = 8'h00;
            12'b01100_1001010: DATA = 8'h00;
            12'b01100_1001011: DATA = 8'h00;
            12'b01100_1001100: DATA = 8'h00;
            12'b01100_1001101: DATA = 8'h00;
            12'b01100_1001110: DATA = 8'h00;
            12'b01100_1001111: DATA = 8'h00;
            // Row 13
            12'b01101_0000000: DATA = 8'h57;
            12'b01101_0000001: DATA = 8'h41;
            12'b01101_0000010: DATA = 8'h56;
            12'b01101_0000011: DATA = 8'h45;
            12'b01101_0000100: DATA = 8'h46;
            12'b01101_0000101: DATA = 8'h4F;
            12'b01101_0000110: DATA = 8'h52;
            12'b01101_0000111: DATA = 8'h4D;
            12'b01101_0001000: DATA = 8'h00;
            12'b01101_0001001: DATA = 8'h00;
            12'b01101_0001010: DATA = 8'h00;
            12'b01101_0001011: DATA = 8'h00;
            12'b01101_0001100: DATA = 8'h00;
            12'b01101_0001101: DATA = 8'h00;
            12'b01101_0001110: DATA = (WAVE2 == 2'b00) ? 8'h53 : (WAVE2 == 2'b01) ? 8'h53 : (WAVE2 == 2'b10) ? 8'h54 : 8'h53;
            12'b01101_0001111: DATA = (WAVE2 == 2'b00) ? 8'h51 : (WAVE2 == 2'b01) ? 8'h41 : (WAVE2 == 2'b10) ? 8'h52 : 8'h49;
            12'b01101_0010000: DATA = (WAVE2 == 2'b00) ? 8'h55 : (WAVE2 == 2'b01) ? 8'h57 : (WAVE2 == 2'b10) ? 8'h49 : 8'h4E;
            12'b01101_0010001: DATA = (WAVE2 == 2'b00) ? 8'h41 : (WAVE2 == 2'b01) ? 8'h54 : (WAVE2 == 2'b10) ? 8'h41 : 8'h45;
            12'b01101_0010010: DATA = (WAVE2 == 2'b00) ? 8'h52 : (WAVE2 == 2'b01) ? 8'h4F : (WAVE2 == 2'b10) ? 8'h4E : 8'h00;
            12'b01101_0010011: DATA = (WAVE2 == 2'b00) ? 8'h45 : (WAVE2 == 2'b01) ? 8'h4F : (WAVE2 == 2'b10) ? 8'h47 : 8'h00;
            12'b01101_0010100: DATA = (WAVE2 == 2'b00) ? 8'h00 : (WAVE2 == 2'b01) ? 8'h54 : (WAVE2 == 2'b10) ? 8'h4C : 8'h00;
            12'b01101_0010101: DATA = (WAVE2 == 2'b00) ? 8'h00 : (WAVE2 == 2'b01) ? 8'h48 : (WAVE2 == 2'b10) ? 8'h45 : 8'h00;
            12'b01101_0010110: DATA = 8'h00;
            12'b01101_0010111: DATA = 8'h00;
            12'b01101_0011000: DATA = 8'h00;
            12'b01101_0011001: DATA = 8'h00;
            12'b01101_0011010: DATA = 8'h00;
            12'b01101_0011011: DATA = 8'h00;
            12'b01101_0011100: DATA = 8'hC6;
            12'b01101_0011101: DATA = (FORM2 == 2'b10 && WAVE2 == 2'b00) ? 8'hA3 : (FORM2 == 2'b10 && WAVE2 == 2'b01) ? 8'hE7 : (FORM2 == 2'b10 && WAVE2 == 2'b10) ? 8'hB7 : (FORM2 == 2'b10 && WAVE2 == 2'b11) ? 8'h8F : 8'h00;
            12'b01101_0011110: DATA = (FORM2 == 2'b10 && WAVE2 == 2'b00) ? 8'hA4 : (FORM2 == 2'b10 && WAVE2 == 2'b01) ? 8'hE8 : (FORM2 == 2'b10 && WAVE2 == 2'b10) ? 8'hB8 : (FORM2 == 2'b10 && WAVE2 == 2'b11) ? 8'h90 : 8'h00;
            12'b01101_0011111: DATA = (FORM2 == 2'b10 && WAVE2 == 2'b00) ? 8'hA5 : (FORM2 == 2'b10 && WAVE2 == 2'b01) ? 8'hE9 : (FORM2 == 2'b10 && WAVE2 == 2'b10) ? 8'hB9 : (FORM2 == 2'b10 && WAVE2 == 2'b11) ? 8'h91 : 8'h00;
            12'b01101_0100000: DATA = (FORM2 == 2'b10 && WAVE2 == 2'b00) ? 8'hA6 : (FORM2 == 2'b10 && WAVE2 == 2'b01) ? 8'hEA : (FORM2 == 2'b10 && WAVE2 == 2'b10) ? 8'hBA : (FORM2 == 2'b10 && WAVE2 == 2'b11) ? 8'h92 : 8'h00;
            12'b01101_0100001: DATA = (FORM2 == 2'b10 && WAVE2 == 2'b00) ? 8'hA7 : (FORM2 == 2'b10 && WAVE2 == 2'b01) ? 8'hEB : (FORM2 == 2'b10 && WAVE2 == 2'b10) ? 8'hBB : (FORM2 == 2'b10 && WAVE2 == 2'b11) ? 8'h93 : 8'h00;
            12'b01101_0100010: DATA = (FORM2 == 2'b01) ? 8'h00 : (FORM2 == 2'b00 && WAVE2 == 2'b00) ? 8'hA3 : (FORM2 == 2'b00 && WAVE2 == 2'b01) ? 8'hCF : (FORM2 == 2'b00 && WAVE2 == 2'b10) ? 8'hB7 : (FORM2 == 2'b00 && WAVE2 == 2'b11) ? 8'h8F : 8'h00;
            12'b01101_0100011: DATA = (FORM2 == 2'b01) ? 8'h00 : (FORM2 == 2'b00 && WAVE2 == 2'b00) ? 8'hA4 : (FORM2 == 2'b00 && WAVE2 == 2'b01) ? 8'hD0 : (FORM2 == 2'b00 && WAVE2 == 2'b10) ? 8'hB8 : (FORM2 == 2'b00 && WAVE2 == 2'b11) ? 8'h90 : 8'h00;
            12'b01101_0100100: DATA = (FORM2 == 2'b01) ? 8'h00 : (FORM2 == 2'b00 && WAVE2 == 2'b00) ? 8'hA5 : (FORM2 == 2'b00 && WAVE2 == 2'b01) ? 8'hD1 : (FORM2 == 2'b00 && WAVE2 == 2'b10) ? 8'hB9 : (FORM2 == 2'b00 && WAVE2 == 2'b11) ? 8'h91 : 8'h00;
            12'b01101_0100101: DATA = (FORM2 == 2'b01) ? 8'h00 : (FORM2 == 2'b00 && WAVE2 == 2'b00) ? 8'hA6 : (FORM2 == 2'b00 && WAVE2 == 2'b01) ? 8'hD2 : (FORM2 == 2'b00 && WAVE2 == 2'b10) ? 8'hBA : (FORM2 == 2'b00 && WAVE2 == 2'b11) ? 8'h92 : 8'h00;
            12'b01101_0100110: DATA = (FORM2 == 2'b01) ? 8'h00 : (FORM2 == 2'b00 && WAVE2 == 2'b00) ? 8'hA7 : (FORM2 == 2'b00 && WAVE2 == 2'b01) ? 8'hD3 : (FORM2 == 2'b00 && WAVE2 == 2'b10) ? 8'hBB : (FORM2 == 2'b00 && WAVE2 == 2'b11) ? 8'h93 : 8'h00;
            12'b01101_0100111: DATA = 8'hC7;
            12'b01101_0101000: DATA = 8'h00;
            12'b01101_0101001: DATA = 8'h00;
            12'b01101_0101010: DATA = 8'h00;
            12'b01101_0101011: DATA = 8'h00;
            12'b01101_0101100: DATA = 8'h00;
            12'b01101_0101101: DATA = 8'h00;
            12'b01101_0101110: DATA = 8'h00;
            12'b01101_0101111: DATA = 8'h00;
            12'b01101_0110000: DATA = 8'h00;
            12'b01101_0110001: DATA = 8'h00;
            12'b01101_0110010: DATA = 8'h00;
            12'b01101_0110011: DATA = 8'h00;
            12'b01101_0110100: DATA = 8'h00;
            12'b01101_0110101: DATA = 8'h00;
            12'b01101_0110110: DATA = 8'h00;
            12'b01101_0110111: DATA = 8'h00;
            12'b01101_0111000: DATA = 8'h00;
            12'b01101_0111001: DATA = 8'h00;
            12'b01101_0111010: DATA = 8'h00;
            12'b01101_0111011: DATA = 8'h00;
            12'b01101_0111100: DATA = 8'h00;
            12'b01101_0111101: DATA = 8'h00;
            12'b01101_0111110: DATA = 8'h00;
            12'b01101_0111111: DATA = 8'h00;
            12'b01101_1000000: DATA = 8'h00;
            12'b01101_1000001: DATA = 8'h00;
            12'b01101_1000010: DATA = 8'h00;
            12'b01101_1000011: DATA = 8'h00;
            12'b01101_1000100: DATA = 8'h00;
            12'b01101_1000101: DATA = 8'h00;
            12'b01101_1000110: DATA = 8'h00;
            12'b01101_1000111: DATA = 8'h00;
            12'b01101_1001000: DATA = 8'h00;
            12'b01101_1001001: DATA = 8'h00;
            12'b01101_1001010: DATA = 8'h00;
            12'b01101_1001011: DATA = 8'h00;
            12'b01101_1001100: DATA = 8'h00;
            12'b01101_1001101: DATA = 8'h00;
            12'b01101_1001110: DATA = 8'h00;
            12'b01101_1001111: DATA = 8'h00;
            // Row 14
            12'b01110_0000000: DATA = 8'h4D;
            12'b01110_0000001: DATA = 8'h4F;
            12'b01110_0000010: DATA = 8'h44;
            12'b01110_0000011: DATA = 8'h45;
            12'b01110_0000100: DATA = 8'h00;
            12'b01110_0000101: DATA = 8'h00;
            12'b01110_0000110: DATA = 8'h00;
            12'b01110_0000111: DATA = 8'h00;
            12'b01110_0001000: DATA = 8'h00;
            12'b01110_0001001: DATA = 8'h00;
            12'b01110_0001010: DATA = 8'h00;
            12'b01110_0001011: DATA = 8'h00;
            12'b01110_0001100: DATA = 8'h00;
            12'b01110_0001101: DATA = 8'h00;
            12'b01110_0001110: DATA = (FORM2 == 2'b00) ? 8'h4E : (FORM2 == 2'b01) ? 8'h48 : (FORM2 == 2'b10) ? 8'h52 : 8'h46;
            12'b01110_0001111: DATA = (FORM2 == 2'b00) ? 8'h4F : (FORM2 == 2'b01) ? 8'h41 : (FORM2 == 2'b10) ? 8'h45 : 8'h55;
            12'b01110_0010000: DATA = (FORM2 == 2'b00) ? 8'h52 : (FORM2 == 2'b01) ? 8'h4C : (FORM2 == 2'b10) ? 8'h56 : 8'h4C;
            12'b01110_0010001: DATA = (FORM2 == 2'b00) ? 8'h4D : (FORM2 == 2'b01) ? 8'h46 : (FORM2 == 2'b10) ? 8'h45 : 8'h4C;
            12'b01110_0010010: DATA = (FORM2 == 2'b00) ? 8'h41 : (FORM2 == 2'b01) ? 8'h2D : (FORM2 == 2'b10) ? 8'h52 : 8'h2D;
            12'b01110_0010011: DATA = (FORM2 == 2'b00) ? 8'h4C : (FORM2 == 2'b01) ? 8'h57 : (FORM2 == 2'b10) ? 8'h53 : 8'h57;
            12'b01110_0010100: DATA = (FORM2 == 2'b00) ? 8'h00 : (FORM2 == 2'b01) ? 8'h41 : (FORM2 == 2'b10) ? 8'h45 : 8'h41;
            12'b01110_0010101: DATA = (FORM2 == 2'b00) ? 8'h00 : (FORM2 == 2'b01) ? 8'h56 : (FORM2 == 2'b10) ? 8'h44 : 8'h56;
            12'b01110_0010110: DATA = (FORM2 == 2'b00) ? 8'h00 : (FORM2 == 2'b01) ? 8'h45 : (FORM2 == 2'b10) ? 8'h00 : 8'h45;
            12'b01110_0010111: DATA = 8'h00;
            12'b01110_0011000: DATA = 8'h00;
            12'b01110_0011001: DATA = 8'h00;
            12'b01110_0011010: DATA = 8'h00;
            12'b01110_0011011: DATA = 8'h00;
            12'b01110_0011100: DATA = 8'hD6;
            12'b01110_0011101: DATA = 8'hC9;
            12'b01110_0011110: DATA = 8'hC9;
            12'b01110_0011111: DATA = 8'hC9;
            12'b01110_0100000: DATA = 8'hC9;
            12'b01110_0100001: DATA = 8'hC9;
            12'b01110_0100010: DATA = 8'hC9;
            12'b01110_0100011: DATA = 8'hC9;
            12'b01110_0100100: DATA = 8'hC9;
            12'b01110_0100101: DATA = 8'hC9;
            12'b01110_0100110: DATA = 8'hC9;
            12'b01110_0100111: DATA = 8'hD7;
            12'b01110_0101000: DATA = 8'h00;
            12'b01110_0101001: DATA = 8'h00;
            12'b01110_0101010: DATA = 8'h00;
            12'b01110_0101011: DATA = 8'h00;
            12'b01110_0101100: DATA = 8'h00;
            12'b01110_0101101: DATA = 8'h00;
            12'b01110_0101110: DATA = 8'h00;
            12'b01110_0101111: DATA = 8'h00;
            12'b01110_0110000: DATA = 8'h00;
            12'b01110_0110001: DATA = 8'h00;
            12'b01110_0110010: DATA = 8'h00;
            12'b01110_0110011: DATA = 8'h00;
            12'b01110_0110100: DATA = 8'h00;
            12'b01110_0110101: DATA = 8'h00;
            12'b01110_0110110: DATA = 8'h00;
            12'b01110_0110111: DATA = 8'h00;
            12'b01110_0111000: DATA = 8'h00;
            12'b01110_0111001: DATA = 8'h00;
            12'b01110_0111010: DATA = 8'h00;
            12'b01110_0111011: DATA = 8'h00;
            12'b01110_0111100: DATA = 8'h00;
            12'b01110_0111101: DATA = 8'h00;
            12'b01110_0111110: DATA = 8'h00;
            12'b01110_0111111: DATA = 8'h00;
            12'b01110_1000000: DATA = 8'h00;
            12'b01110_1000001: DATA = 8'h00;
            12'b01110_1000010: DATA = 8'h00;
            12'b01110_1000011: DATA = 8'h00;
            12'b01110_1000100: DATA = 8'h00;
            12'b01110_1000101: DATA = 8'h00;
            12'b01110_1000110: DATA = 8'h00;
            12'b01110_1000111: DATA = 8'h00;
            12'b01110_1001000: DATA = 8'h00;
            12'b01110_1001001: DATA = 8'h00;
            12'b01110_1001010: DATA = 8'h00;
            12'b01110_1001011: DATA = 8'h00;
            12'b01110_1001100: DATA = 8'h00;
            12'b01110_1001101: DATA = 8'h00;
            12'b01110_1001110: DATA = 8'h00;
            12'b01110_1001111: DATA = 8'h00;
            // Row 15
            12'b01111_0000000: DATA = 8'h00;
            12'b01111_0000001: DATA = 8'h00;
            12'b01111_0000010: DATA = 8'h00;
            12'b01111_0000011: DATA = 8'h00;
            12'b01111_0000100: DATA = 8'h00;
            12'b01111_0000101: DATA = 8'h00;
            12'b01111_0000110: DATA = 8'h00;
            12'b01111_0000111: DATA = 8'h00;
            12'b01111_0001000: DATA = 8'h00;
            12'b01111_0001001: DATA = 8'h00;
            12'b01111_0001010: DATA = 8'h00;
            12'b01111_0001011: DATA = 8'h00;
            12'b01111_0001100: DATA = 8'h00;
            12'b01111_0001101: DATA = 8'h00;
            12'b01111_0001110: DATA = 8'h00;
            12'b01111_0001111: DATA = 8'h00;
            12'b01111_0010000: DATA = 8'h00;
            12'b01111_0010001: DATA = 8'h00;
            12'b01111_0010010: DATA = 8'h00;
            12'b01111_0010011: DATA = 8'h00;
            12'b01111_0010100: DATA = 8'h00;
            12'b01111_0010101: DATA = 8'h00;
            12'b01111_0010110: DATA = 8'h00;
            12'b01111_0010111: DATA = 8'h00;
            12'b01111_0011000: DATA = 8'h00;
            12'b01111_0011001: DATA = 8'h00;
            12'b01111_0011010: DATA = 8'h00;
            12'b01111_0011011: DATA = 8'h00;
            12'b01111_0011100: DATA = 8'h00;
            12'b01111_0011101: DATA = 8'h00;
            12'b01111_0011110: DATA = 8'h00;
            12'b01111_0011111: DATA = 8'h00;
            12'b01111_0100000: DATA = 8'h00;
            12'b01111_0100001: DATA = 8'h00;
            12'b01111_0100010: DATA = 8'h00;
            12'b01111_0100011: DATA = 8'h00;
            12'b01111_0100100: DATA = 8'h00;
            12'b01111_0100101: DATA = 8'h00;
            12'b01111_0100110: DATA = 8'h00;
            12'b01111_0100111: DATA = 8'h00;
            12'b01111_0101000: DATA = 8'h00;
            12'b01111_0101001: DATA = 8'h00;
            12'b01111_0101010: DATA = 8'h00;
            12'b01111_0101011: DATA = 8'h00;
            12'b01111_0101100: DATA = 8'h00;
            12'b01111_0101101: DATA = 8'h00;
            12'b01111_0101110: DATA = 8'h00;
            12'b01111_0101111: DATA = 8'h00;
            12'b01111_0110000: DATA = 8'h00;
            12'b01111_0110001: DATA = 8'h00;
            12'b01111_0110010: DATA = 8'h00;
            12'b01111_0110011: DATA = 8'h00;
            12'b01111_0110100: DATA = 8'h00;
            12'b01111_0110101: DATA = 8'h00;
            12'b01111_0110110: DATA = 8'h00;
            12'b01111_0110111: DATA = 8'h00;
            12'b01111_0111000: DATA = 8'h00;
            12'b01111_0111001: DATA = 8'h00;
            12'b01111_0111010: DATA = 8'h00;
            12'b01111_0111011: DATA = 8'h00;
            12'b01111_0111100: DATA = 8'h00;
            12'b01111_0111101: DATA = 8'h00;
            12'b01111_0111110: DATA = 8'h00;
            12'b01111_0111111: DATA = 8'h00;
            12'b01111_1000000: DATA = 8'h00;
            12'b01111_1000001: DATA = 8'h00;
            12'b01111_1000010: DATA = 8'h00;
            12'b01111_1000011: DATA = 8'h00;
            12'b01111_1000100: DATA = 8'h00;
            12'b01111_1000101: DATA = 8'h00;
            12'b01111_1000110: DATA = 8'h00;
            12'b01111_1000111: DATA = 8'h00;
            12'b01111_1001000: DATA = 8'h00;
            12'b01111_1001001: DATA = 8'h00;
            12'b01111_1001010: DATA = 8'h00;
            12'b01111_1001011: DATA = 8'h00;
            12'b01111_1001100: DATA = 8'h00;
            12'b01111_1001101: DATA = 8'h00;
            12'b01111_1001110: DATA = 8'h00;
            12'b01111_1001111: DATA = 8'h00;
            // Row 16
            12'b10000_0000000: DATA = 8'h4D;
            12'b10000_0000001: DATA = 8'h49;
            12'b10000_0000010: DATA = 8'h4E;
            12'b10000_0000011: DATA = 8'h00;
            12'b10000_0000100: DATA = (WAVE == 1) ? 8'h00 : (MIN_MAX == 0) ? 8'h3C : (BOTH == 1) ? 8'h3C : 8'h00;
            12'b10000_0000101: DATA = 8'h00;
            12'b10000_0000110: DATA = 8'h00;
            12'b10000_0000111: DATA = 8'h00;
            12'b10000_0001000: DATA = 8'h00;
            12'b10000_0001001: DATA = 8'h4D;
            12'b10000_0001010: DATA = 8'h41;
            12'b10000_0001011: DATA = 8'h58;
            12'b10000_0001100: DATA = 8'h00;
            12'b10000_0001101: DATA = (WAVE == 1) ? 8'h00 : (MIN_MAX == 1) ? 8'h3C : (BOTH == 1) ? 8'h3C : 8'h00;
            12'b10000_0001110: DATA = 8'h00;
            12'b10000_0001111: DATA = 8'h00;
            12'b10000_0010000: DATA = 8'h00;
            12'b10000_0010001: DATA = 8'h00;
            12'b10000_0010010: DATA = 8'h00;
            12'b10000_0010011: DATA = 8'h00;
            12'b10000_0010100: DATA = 8'h00;
            12'b10000_0010101: DATA = 8'h00;
            12'b10000_0010110: DATA = 8'h00;
            12'b10000_0010111: DATA = 8'h00;
            12'b10000_0011000: DATA = 8'h00;
            12'b10000_0011001: DATA = 8'h00;
            12'b10000_0011010: DATA = 8'h00;
            12'b10000_0011011: DATA = 8'h00;
            12'b10000_0011100: DATA = (WAVE1 == 2'b00 && CHANNEL == 0 || WAVE1 == 2'b10 && CHANNEL == 0 || WAVE2 == 2'b00 && CHANNEL == 1 || WAVE2 == 2'b10 && CHANNEL == 1) ? 8'h44 : 8'h00;
            12'b10000_0011101: DATA = (WAVE1 == 2'b00 && CHANNEL == 0 || WAVE1 == 2'b10 && CHANNEL == 0 || WAVE2 == 2'b00 && CHANNEL == 1 || WAVE2 == 2'b10 && CHANNEL == 1) ? 8'h55 : 8'h00;
            12'b10000_0011110: DATA = (WAVE1 == 2'b00 && CHANNEL == 0 || WAVE1 == 2'b10 && CHANNEL == 0 || WAVE2 == 2'b00 && CHANNEL == 1 || WAVE2 == 2'b10 && CHANNEL == 1) ? 8'h54 : 8'h00;
            12'b10000_0011111: DATA = (WAVE1 == 2'b00 && CHANNEL == 0 || WAVE1 == 2'b10 && CHANNEL == 0 || WAVE2 == 2'b00 && CHANNEL == 1 || WAVE2 == 2'b10 && CHANNEL == 1) ? 8'h59 : 8'h00;
            12'b10000_0100000: DATA = 8'h00;
            12'b10000_0100001: DATA = (WAVE1 == 2'b00 && CHANNEL == 0 || WAVE1 == 2'b10 && CHANNEL == 0 || WAVE2 == 2'b00 && CHANNEL == 1 || WAVE2 == 2'b10 && CHANNEL == 1) ? 8'h43 : 8'h00;
            12'b10000_0100010: DATA = (WAVE1 == 2'b00 && CHANNEL == 0 || WAVE1 == 2'b10 && CHANNEL == 0 || WAVE2 == 2'b00 && CHANNEL == 1 || WAVE2 == 2'b10 && CHANNEL == 1) ? 8'h59 : 8'h00;
            12'b10000_0100011: DATA = (WAVE1 == 2'b00 && CHANNEL == 0 || WAVE1 == 2'b10 && CHANNEL == 0 || WAVE2 == 2'b00 && CHANNEL == 1 || WAVE2 == 2'b10 && CHANNEL == 1) ? 8'h43 : 8'h00;
            12'b10000_0100100: DATA = (WAVE1 == 2'b00 && CHANNEL == 0 || WAVE1 == 2'b10 && CHANNEL == 0 || WAVE2 == 2'b00 && CHANNEL == 1 || WAVE2 == 2'b10 && CHANNEL == 1) ? 8'h4C : 8'h00;
            12'b10000_0100101: DATA = (WAVE1 == 2'b00 && CHANNEL == 0 || WAVE1 == 2'b10 && CHANNEL == 0 || WAVE2 == 2'b00 && CHANNEL == 1 || WAVE2 == 2'b10 && CHANNEL == 1) ? 8'h45 : 8'h00;
            12'b10000_0100110: DATA = 8'h00;
            12'b10000_0100111: DATA = (WAVE1 == 2'b00 && CHANNEL == 0 || WAVE1 == 2'b10 && CHANNEL == 0 || WAVE2 == 2'b00 && CHANNEL == 1 || WAVE2 == 2'b10 && CHANNEL == 1) ? DUTY_CYCLE[23:16] : 8'h00;
            12'b10000_0101000: DATA = (WAVE1 == 2'b00 && CHANNEL == 0 || WAVE1 == 2'b10 && CHANNEL == 0 || WAVE2 == 2'b00 && CHANNEL == 1 || WAVE2 == 2'b10 && CHANNEL == 1) ? DUTY_CYCLE[15:8] : 8'h00;
            12'b10000_0101001: DATA = (WAVE1 == 2'b00 && CHANNEL == 0 || WAVE1 == 2'b10 && CHANNEL == 0 || WAVE2 == 2'b00 && CHANNEL == 1 || WAVE2 == 2'b10 && CHANNEL == 1) ? DUTY_CYCLE[7:0] : 8'h00;
            12'b10000_0101010: DATA = 8'h00;
            12'b10000_0101011: DATA = 8'h00;
            12'b10000_0101100: DATA = 8'h00;
            12'b10000_0101101: DATA = 8'h00;
            12'b10000_0101110: DATA = 8'h00;
            12'b10000_0101111: DATA = 8'h00;
            12'b10000_0110000: DATA = 8'h00;
            12'b10000_0110001: DATA = 8'h00;
            12'b10000_0110010: DATA = 8'h00;
            12'b10000_0110011: DATA = 8'h00;
            12'b10000_0110100: DATA = 8'h00;
            12'b10000_0110101: DATA = 8'h00;
            12'b10000_0110110: DATA = 8'h00;
            12'b10000_0110111: DATA = 8'h00;
            12'b10000_0111000: DATA = 8'h00;
            12'b10000_0111001: DATA = 8'h00;
            12'b10000_0111010: DATA = 8'h00;
            12'b10000_0111011: DATA = 8'h00;
            12'b10000_0111100: DATA = 8'h00;
            12'b10000_0111101: DATA = 8'h00;
            12'b10000_0111110: DATA = 8'h00;
            12'b10000_0111111: DATA = 8'h00;
            12'b10000_1000000: DATA = 8'h00;
            12'b10000_1000001: DATA = 8'h00;
            12'b10000_1000010: DATA = 8'h00;
            12'b10000_1000011: DATA = 8'h00;
            12'b10000_1000100: DATA = 8'h00;
            12'b10000_1000101: DATA = 8'h00;
            12'b10000_1000110: DATA = 8'h00;
            12'b10000_1000111: DATA = 8'h00;
            12'b10000_1001000: DATA = 8'h00;
            12'b10000_1001001: DATA = 8'h00;
            12'b10000_1001010: DATA = 8'h00;
            12'b10000_1001011: DATA = 8'h00;
            12'b10000_1001100: DATA = 8'h00;
            12'b10000_1001101: DATA = 8'h00;
            12'b10000_1001110: DATA = 8'h00;
            12'b10000_1001111: DATA = 8'h00;
            // Row 17
            12'b10001_0000000: DATA = 8'h43;
            12'b10001_0000001: DATA = 8'h48;
            12'b10001_0000010: DATA = 8'h41;
            12'b10001_0000011: DATA = 8'h4E;
            12'b10001_0000100: DATA = 8'h47;
            12'b10001_0000101: DATA = 8'h45;
            12'b10001_0000110: DATA = 8'h00;
            12'b10001_0000111: DATA = 8'h57;
            12'b10001_0001000: DATA = 8'h41;
            12'b10001_0001001: DATA = 8'h56;
            12'b10001_0001010: DATA = 8'h45;
            12'b10001_0001011: DATA = 8'h00;
            12'b10001_0001100: DATA = 8'h00;
            12'b10001_0001101: DATA = 8'h00;
            12'b10001_0001110: DATA = 8'h4F;
            12'b10001_0001111: DATA = (WAVE == 1) ? 8'h4E : 8'h46;
            12'b10001_0010000: DATA = (WAVE == 1) ? 8'h00 : 8'h46;
            12'b10001_0010001: DATA = 8'h00;
            12'b10001_0010010: DATA = 8'h00;
            12'b10001_0010011: DATA = 8'h00;
            12'b10001_0010100: DATA = 8'h00;
            12'b10001_0010101: DATA = 8'h00;
            12'b10001_0010110: DATA = 8'h00;
            12'b10001_0010111: DATA = 8'h00;
            12'b10001_0011000: DATA = 8'h00;
            12'b10001_0011001: DATA = 8'h00;
            12'b10001_0011010: DATA = 8'h00;
            12'b10001_0011011: DATA = 8'h00;
            12'b10001_0011100: DATA = 8'h00;
            12'b10001_0011101: DATA = 8'h00;
            12'b10001_0011110: DATA = 8'h00;
            12'b10001_0011111: DATA = 8'h00;
            12'b10001_0100000: DATA = 8'h00;
            12'b10001_0100001: DATA = 8'h00;
            12'b10001_0100010: DATA = 8'h00;
            12'b10001_0100011: DATA = 8'h00;
            12'b10001_0100100: DATA = 8'h00;
            12'b10001_0100101: DATA = 8'h00;
            12'b10001_0100110: DATA = 8'h00;
            12'b10001_0100111: DATA = 8'h00;
            12'b10001_0101000: DATA = 8'h00;
            12'b10001_0101001: DATA = 8'h00;
            12'b10001_0101010: DATA = 8'h00;
            12'b10001_0101011: DATA = 8'h00;
            12'b10001_0101100: DATA = 8'h00;
            12'b10001_0101101: DATA = 8'h00;
            12'b10001_0101110: DATA = 8'h00;
            12'b10001_0101111: DATA = 8'h00;
            12'b10001_0110000: DATA = 8'h00;
            12'b10001_0110001: DATA = 8'h00;
            12'b10001_0110010: DATA = 8'h00;
            12'b10001_0110011: DATA = 8'h00;
            12'b10001_0110100: DATA = 8'h00;
            12'b10001_0110101: DATA = 8'h00;
            12'b10001_0110110: DATA = 8'h00;
            12'b10001_0110111: DATA = 8'h00;
            12'b10001_0111000: DATA = 8'h00;
            12'b10001_0111001: DATA = 8'h00;
            12'b10001_0111010: DATA = 8'h00;
            12'b10001_0111011: DATA = 8'h00;
            12'b10001_0111100: DATA = 8'h00;
            12'b10001_0111101: DATA = 8'h00;
            12'b10001_0111110: DATA = 8'h00;
            12'b10001_0111111: DATA = 8'h00;
            12'b10001_1000000: DATA = 8'h00;
            12'b10001_1000001: DATA = 8'h00;
            12'b10001_1000010: DATA = 8'h00;
            12'b10001_1000011: DATA = 8'h00;
            12'b10001_1000100: DATA = 8'h00;
            12'b10001_1000101: DATA = 8'h00;
            12'b10001_1000110: DATA = 8'h00;
            12'b10001_1000111: DATA = 8'h00;
            12'b10001_1001000: DATA = 8'h00;
            12'b10001_1001001: DATA = 8'h00;
            12'b10001_1001010: DATA = 8'h00;
            12'b10001_1001011: DATA = 8'h00;
            12'b10001_1001100: DATA = 8'h00;
            12'b10001_1001101: DATA = 8'h00;
            12'b10001_1001110: DATA = 8'h00;
            12'b10001_1001111: DATA = 8'h00;
            // Row 18
            12'b10010_0000000: DATA = 8'h4B;
            12'b10010_0000001: DATA = 8'h45;
            12'b10010_0000010: DATA = 8'h59;
            12'b10010_0000011: DATA = 8'h42;
            12'b10010_0000100: DATA = 8'h4F;
            12'b10010_0000101: DATA = 8'h41;
            12'b10010_0000110: DATA = 8'h52;
            12'b10010_0000111: DATA = 8'h44;
            12'b10010_0001000: DATA = 8'h00;
            12'b10010_0001001: DATA = 8'h00;
            12'b10010_0001010: DATA = 8'h00;
            12'b10010_0001011: DATA = 8'h00;
            12'b10010_0001100: DATA = 8'h00;
            12'b10010_0001101: DATA = 8'h00;
            12'b10010_0001110: DATA = 8'h4F;
            12'b10010_0001111: DATA = (KEYBOARD == 1) ? 8'h4E : 8'h46;
            12'b10010_0010000: DATA = (KEYBOARD == 1) ? 8'h00 : 8'h46;
            12'b10010_0010001: DATA = 8'h00;
            12'b10010_0010010: DATA = 8'h00;
            12'b10010_0010011: DATA = 8'h00;
            12'b10010_0010100: DATA = 8'h00;
            12'b10010_0010101: DATA = 8'h00;
            12'b10010_0010110: DATA = 8'h00;
            12'b10010_0010111: DATA = 8'h00;
            12'b10010_0011000: DATA = 8'h00;
            12'b10010_0011001: DATA = 8'h00;
            12'b10010_0011010: DATA = 8'h00;
            12'b10010_0011011: DATA = 8'h00;
            12'b10010_0011100: DATA = 8'h00;
            12'b10010_0011101: DATA = 8'h00;
            12'b10010_0011110: DATA = 8'h00;
            12'b10010_0011111: DATA = 8'h00;
            12'b10010_0100000: DATA = 8'h00;
            12'b10010_0100001: DATA = 8'h00;
            12'b10010_0100010: DATA = 8'h00;
            12'b10010_0100011: DATA = 8'h00;
            12'b10010_0100100: DATA = 8'h00;
            12'b10010_0100101: DATA = 8'h00;
            12'b10010_0100110: DATA = 8'h00;
            12'b10010_0100111: DATA = 8'h00;
            12'b10010_0101000: DATA = 8'h00;
            12'b10010_0101001: DATA = 8'h00;
            12'b10010_0101010: DATA = 8'h00;
            12'b10010_0101011: DATA = 8'h00;
            12'b10010_0101100: DATA = 8'h00;
            12'b10010_0101101: DATA = 8'h00;
            12'b10010_0101110: DATA = 8'h00;
            12'b10010_0101111: DATA = 8'h00;
            12'b10010_0110000: DATA = 8'h00;
            12'b10010_0110001: DATA = 8'h00;
            12'b10010_0110010: DATA = 8'h00;
            12'b10010_0110011: DATA = 8'h00;
            12'b10010_0110100: DATA = 8'h00;
            12'b10010_0110101: DATA = 8'h00;
            12'b10010_0110110: DATA = 8'h00;
            12'b10010_0110111: DATA = 8'h00;
            12'b10010_0111000: DATA = 8'h00;
            12'b10010_0111001: DATA = 8'h00;
            12'b10010_0111010: DATA = 8'h00;
            12'b10010_0111011: DATA = 8'h00;
            12'b10010_0111100: DATA = 8'h00;
            12'b10010_0111101: DATA = 8'h00;
            12'b10010_0111110: DATA = 8'h00;
            12'b10010_0111111: DATA = 8'h00;
            12'b10010_1000000: DATA = 8'h00;
            12'b10010_1000001: DATA = 8'h00;
            12'b10010_1000010: DATA = 8'h00;
            12'b10010_1000011: DATA = 8'h00;
            12'b10010_1000100: DATA = 8'h00;
            12'b10010_1000101: DATA = 8'h00;
            12'b10010_1000110: DATA = 8'h00;
            12'b10010_1000111: DATA = 8'h00;
            12'b10010_1001000: DATA = 8'h00;
            12'b10010_1001001: DATA = 8'h00;
            12'b10010_1001010: DATA = 8'h00;
            12'b10010_1001011: DATA = 8'h00;
            12'b10010_1001100: DATA = 8'h00;
            12'b10010_1001101: DATA = 8'h00;
            12'b10010_1001110: DATA = 8'h00;
            12'b10010_1001111: DATA = 8'h00;
            // Row 19
            12'b10011_0000000: DATA = 8'h4D;
            12'b10011_0000001: DATA = 8'h41;
            12'b10011_0000010: DATA = 8'h58;
            12'b10011_0000011: DATA = 8'h00;
            12'b10011_0000100: DATA = 8'h41;
            12'b10011_0000101: DATA = 8'h4D;
            12'b10011_0000110: DATA = 8'h50;
            12'b10011_0000111: DATA = 8'h00;
            12'b10011_0001000: DATA = 8'h4D;
            12'b10011_0001001: DATA = 8'h4F;
            12'b10011_0001010: DATA = 8'h44;
            12'b10011_0001011: DATA = 8'h00;
            12'b10011_0001100: DATA = 8'h00;
            12'b10011_0001101: DATA = 8'h00;
            12'b10011_0001110: DATA = 8'h4F;
            12'b10011_0001111: DATA = (MAX_AMP_MOD == 1) ? 8'h4E : 8'h46;
            12'b10011_0010000: DATA = (MAX_AMP_MOD == 1) ? 8'h00 : 8'h46;
            12'b10011_0010001: DATA = 8'h00;
            12'b10011_0010010: DATA = 8'h00;
            12'b10011_0010011: DATA = 8'h00;
            12'b10011_0010100: DATA = 8'h00;
            12'b10011_0010101: DATA = 8'h00;
            12'b10011_0010110: DATA = 8'h00;
            12'b10011_0010111: DATA = 8'h00;
            12'b10011_0011000: DATA = 8'h00;
            12'b10011_0011001: DATA = 8'h00;
            12'b10011_0011010: DATA = 8'h00;
            12'b10011_0011011: DATA = 8'h00;
            12'b10011_0011100: DATA = 8'h00;
            12'b10011_0011101: DATA = 8'h00;
            12'b10011_0011110: DATA = 8'h00;
            12'b10011_0011111: DATA = 8'h00;
            12'b10011_0100000: DATA = 8'h00;
            12'b10011_0100001: DATA = 8'h00;
            12'b10011_0100010: DATA = 8'h00;
            12'b10011_0100011: DATA = 8'h00;
            12'b10011_0100100: DATA = 8'h00;
            12'b10011_0100101: DATA = 8'h00;
            12'b10011_0100110: DATA = 8'h00;
            12'b10011_0100111: DATA = 8'h00;
            12'b10011_0101000: DATA = 8'h00;
            12'b10011_0101001: DATA = 8'h00;
            12'b10011_0101010: DATA = 8'h00;
            12'b10011_0101011: DATA = 8'h00;
            12'b10011_0101100: DATA = 8'h00;
            12'b10011_0101101: DATA = 8'h00;
            12'b10011_0101110: DATA = 8'h00;
            12'b10011_0101111: DATA = 8'h00;
            12'b10011_0110000: DATA = 8'h00;
            12'b10011_0110001: DATA = 8'h00;
            12'b10011_0110010: DATA = 8'h00;
            12'b10011_0110011: DATA = 8'h00;
            12'b10011_0110100: DATA = 8'h00;
            12'b10011_0110101: DATA = 8'h00;
            12'b10011_0110110: DATA = 8'h00;
            12'b10011_0110111: DATA = 8'h00;
            12'b10011_0111000: DATA = 8'h00;
            12'b10011_0111001: DATA = 8'h00;
            12'b10011_0111010: DATA = 8'h00;
            12'b10011_0111011: DATA = 8'h00;
            12'b10011_0111100: DATA = 8'h00;
            12'b10011_0111101: DATA = 8'h00;
            12'b10011_0111110: DATA = 8'h00;
            12'b10011_0111111: DATA = 8'h00;
            12'b10011_1000000: DATA = 8'h00;
            12'b10011_1000001: DATA = 8'h00;
            12'b10011_1000010: DATA = 8'h00;
            12'b10011_1000011: DATA = 8'h00;
            12'b10011_1000100: DATA = 8'h00;
            12'b10011_1000101: DATA = 8'h00;
            12'b10011_1000110: DATA = 8'h00;
            12'b10011_1000111: DATA = 8'h00;
            12'b10011_1001000: DATA = 8'h00;
            12'b10011_1001001: DATA = 8'h00;
            12'b10011_1001010: DATA = 8'h00;
            12'b10011_1001011: DATA = 8'h00;
            12'b10011_1001100: DATA = 8'h00;
            12'b10011_1001101: DATA = 8'h00;
            12'b10011_1001110: DATA = 8'h00;
            12'b10011_1001111: DATA = 8'h00;
            // Row 20
            12'b10100_0000000: DATA = 8'h4D;
            12'b10100_0000001: DATA = 8'h49;
            12'b10100_0000010: DATA = 8'h4E;
            12'b10100_0000011: DATA = 8'h00;
            12'b10100_0000100: DATA = 8'h4D;
            12'b10100_0000101: DATA = 8'h41;
            12'b10100_0000110: DATA = 8'h58;
            12'b10100_0000111: DATA = 8'h00;
            12'b10100_0001000: DATA = 8'h4D;
            12'b10100_0001001: DATA = 8'h4F;
            12'b10100_0001010: DATA = 8'h44;
            12'b10100_0001011: DATA = 8'h00;
            12'b10100_0001100: DATA = 8'h00;
            12'b10100_0001101: DATA = 8'h00;
            12'b10100_0001110: DATA = 8'h4F;
            12'b10100_0001111: DATA = (MIN_MAX_AMP_MOD == 1) ? 8'h4E : 8'h46;
            12'b10100_0010000: DATA = (MIN_MAX_AMP_MOD == 1) ? 8'h00 : 8'h46;
            12'b10100_0010001: DATA = 8'h00;
            12'b10100_0010010: DATA = 8'h00;
            12'b10100_0010011: DATA = 8'h00;
            12'b10100_0010100: DATA = 8'h00;
            12'b10100_0010101: DATA = 8'h00;
            12'b10100_0010110: DATA = 8'h00;
            12'b10100_0010111: DATA = 8'h00;
            12'b10100_0011000: DATA = 8'h00;
            12'b10100_0011001: DATA = 8'h00;
            12'b10100_0011010: DATA = 8'h00;
            12'b10100_0011011: DATA = 8'h00;
            12'b10100_0011100: DATA = 8'h00;
            12'b10100_0011101: DATA = 8'h00;
            12'b10100_0011110: DATA = 8'h00;
            12'b10100_0011111: DATA = 8'h00;
            12'b10100_0100000: DATA = 8'h00;
            12'b10100_0100001: DATA = 8'h00;
            12'b10100_0100010: DATA = 8'h00;
            12'b10100_0100011: DATA = 8'h00;
            12'b10100_0100100: DATA = 8'h00;
            12'b10100_0100101: DATA = 8'h00;
            12'b10100_0100110: DATA = 8'h00;
            12'b10100_0100111: DATA = 8'h00;
            12'b10100_0101000: DATA = 8'h00;
            12'b10100_0101001: DATA = 8'h00;
            12'b10100_0101010: DATA = 8'h00;
            12'b10100_0101011: DATA = 8'h00;
            12'b10100_0101100: DATA = 8'h00;
            12'b10100_0101101: DATA = 8'h00;
            12'b10100_0101110: DATA = 8'h00;
            12'b10100_0101111: DATA = 8'h00;
            12'b10100_0110000: DATA = 8'h00;
            12'b10100_0110001: DATA = 8'h00;
            12'b10100_0110010: DATA = 8'h00;
            12'b10100_0110011: DATA = 8'h00;
            12'b10100_0110100: DATA = 8'h00;
            12'b10100_0110101: DATA = 8'h00;
            12'b10100_0110110: DATA = 8'h00;
            12'b10100_0110111: DATA = 8'h00;
            12'b10100_0111000: DATA = 8'h00;
            12'b10100_0111001: DATA = 8'h00;
            12'b10100_0111010: DATA = 8'h00;
            12'b10100_0111011: DATA = 8'h00;
            12'b10100_0111100: DATA = 8'h00;
            12'b10100_0111101: DATA = 8'h00;
            12'b10100_0111110: DATA = 8'h00;
            12'b10100_0111111: DATA = 8'h00;
            12'b10100_1000000: DATA = 8'h00;
            12'b10100_1000001: DATA = 8'h00;
            12'b10100_1000010: DATA = 8'h00;
            12'b10100_1000011: DATA = 8'h00;
            12'b10100_1000100: DATA = 8'h00;
            12'b10100_1000101: DATA = 8'h00;
            12'b10100_1000110: DATA = 8'h00;
            12'b10100_1000111: DATA = 8'h00;
            12'b10100_1001000: DATA = 8'h00;
            12'b10100_1001001: DATA = 8'h00;
            12'b10100_1001010: DATA = 8'h00;
            12'b10100_1001011: DATA = 8'h00;
            12'b10100_1001100: DATA = 8'h00;
            12'b10100_1001101: DATA = 8'h00;
            12'b10100_1001110: DATA = 8'h00;
            12'b10100_1001111: DATA = 8'h00;
            // Row 21
            12'b10101_0000000: DATA = 8'h46;
            12'b10101_0000001: DATA = 8'h52;
            12'b10101_0000010: DATA = 8'h45;
            12'b10101_0000011: DATA = 8'h51;
            12'b10101_0000100: DATA = 8'h00;
            12'b10101_0000101: DATA = 8'h4D;
            12'b10101_0000110: DATA = 8'h4F;
            12'b10101_0000111: DATA = 8'h44;
            12'b10101_0001000: DATA = 8'h00;
            12'b10101_0001001: DATA = 8'h00;
            12'b10101_0001010: DATA = 8'h00;
            12'b10101_0001011: DATA = 8'h00;
            12'b10101_0001100: DATA = 8'h00;
            12'b10101_0001101: DATA = 8'h00;
            12'b10101_0001110: DATA = 8'h4F;
            12'b10101_0001111: DATA = (FREQ_MOD == 1) ? 8'h4E : 8'h46;
            12'b10101_0010000: DATA = (FREQ_MOD == 1) ? 8'h00 : 8'h46;
            12'b10101_0010001: DATA = 8'h00;
            12'b10101_0010010: DATA = 8'h00;
            12'b10101_0010011: DATA = 8'h00;
            12'b10101_0010100: DATA = 8'h00;
            12'b10101_0010101: DATA = 8'h00;
            12'b10101_0010110: DATA = 8'h00;
            12'b10101_0010111: DATA = 8'h00;
            12'b10101_0011000: DATA = 8'h00;
            12'b10101_0011001: DATA = 8'h00;
            12'b10101_0011010: DATA = 8'h00;
            12'b10101_0011011: DATA = 8'h00;
            12'b10101_0011100: DATA = (FREQ_MOD == 1) ? 8'h42 : 8'h00;
            12'b10101_0011101: DATA = (FREQ_MOD == 1) ? 8'h41 : 8'h00;
            12'b10101_0011110: DATA = (FREQ_MOD == 1) ? 8'h4E : 8'h00;
            12'b10101_0011111: DATA = (FREQ_MOD == 1) ? 8'h44 : 8'h00;
            12'b10101_0100000: DATA = (FREQ_MOD == 1) ? 8'h57 : 8'h00;
            12'b10101_0100001: DATA = (FREQ_MOD == 1) ? 8'h49 : 8'h00;
            12'b10101_0100010: DATA = (FREQ_MOD == 1) ? 8'h44 : 8'h00;
            12'b10101_0100011: DATA = (FREQ_MOD == 1) ? 8'h54 : 8'h00;
            12'b10101_0100100: DATA = (FREQ_MOD == 1) ? 8'h48 : 8'h00;
            12'b10101_0100101: DATA = 8'h00;
            12'b10101_0100110: DATA = (FREQ_MOD == 1) ? BANDWIDTH[23:16] : 8'h00;
            12'b10101_0100111: DATA = (FREQ_MOD == 1) ? BANDWIDTH[15:8] : 8'h00;
            12'b10101_0101000: DATA = (FREQ_MOD == 1) ? BANDWIDTH[7:0] : 8'h00;
            12'b10101_0101001: DATA = 8'h00;
            12'b10101_0101010: DATA = 8'h00;
            12'b10101_0101011: DATA = 8'h00;
            12'b10101_0101100: DATA = 8'h00;
            12'b10101_0101101: DATA = 8'h00;
            12'b10101_0101110: DATA = 8'h00;
            12'b10101_0101111: DATA = 8'h00;
            12'b10101_0110000: DATA = 8'h00;
            12'b10101_0110001: DATA = 8'h00;
            12'b10101_0110010: DATA = 8'h00;
            12'b10101_0110011: DATA = 8'h00;
            12'b10101_0110100: DATA = 8'h00;
            12'b10101_0110101: DATA = 8'h00;
            12'b10101_0110110: DATA = 8'h00;
            12'b10101_0110111: DATA = 8'h00;
            12'b10101_0111000: DATA = 8'h00;
            12'b10101_0111001: DATA = 8'h00;
            12'b10101_0111010: DATA = 8'h00;
            12'b10101_0111011: DATA = 8'h00;
            12'b10101_0111100: DATA = 8'h00;
            12'b10101_0111101: DATA = 8'h00;
            12'b10101_0111110: DATA = 8'h00;
            12'b10101_0111111: DATA = 8'h00;
            12'b10101_1000000: DATA = 8'h00;
            12'b10101_1000001: DATA = 8'h00;
            12'b10101_1000010: DATA = 8'h00;
            12'b10101_1000011: DATA = 8'h00;
            12'b10101_1000100: DATA = 8'h00;
            12'b10101_1000101: DATA = 8'h00;
            12'b10101_1000110: DATA = 8'h00;
            12'b10101_1000111: DATA = 8'h00;
            12'b10101_1001000: DATA = 8'h00;
            12'b10101_1001001: DATA = 8'h00;
            12'b10101_1001010: DATA = 8'h00;
            12'b10101_1001011: DATA = 8'h00;
            12'b10101_1001100: DATA = 8'h00;
            12'b10101_1001101: DATA = 8'h00;
            12'b10101_1001110: DATA = 8'h00;
            12'b10101_1001111: DATA = 8'h00;
            // Row 22
            12'b10110_0000000: DATA = 8'h50;
            12'b10110_0000001: DATA = 8'h48;
            12'b10110_0000010: DATA = 8'h41;
            12'b10110_0000011: DATA = 8'h53;
            12'b10110_0000100: DATA = 8'h45;
            12'b10110_0000101: DATA = 8'h00;
            12'b10110_0000110: DATA = 8'h4D;
            12'b10110_0000111: DATA = 8'h4F;
            12'b10110_0001000: DATA = 8'h44;
            12'b10110_0001001: DATA = 8'h00;
            12'b10110_0001010: DATA = 8'h00;
            12'b10110_0001011: DATA = 8'h00;
            12'b10110_0001100: DATA = 8'h00;
            12'b10110_0001101: DATA = 8'h00;
            12'b10110_0001110: DATA = 8'h4F;
            12'b10110_0001111: DATA = (PHASE_MOD == 1) ? 8'h4E : 8'h46;
            12'b10110_0010000: DATA = (PHASE_MOD == 1) ? 8'h00 : 8'h46;
            12'b10110_0010001: DATA = 8'h00;
            12'b10110_0010010: DATA = 8'h00;
            12'b10110_0010011: DATA = 8'h00;
            12'b10110_0010100: DATA = 8'h00;
            12'b10110_0010101: DATA = 8'h00;
            12'b10110_0010110: DATA = 8'h00;
            12'b10110_0010111: DATA = 8'h00;
            12'b10110_0011000: DATA = 8'h00;
            12'b10110_0011001: DATA = 8'h00;
            12'b10110_0011010: DATA = 8'h00;
            12'b10110_0011011: DATA = 8'h00;
            12'b10110_0011100: DATA = 8'h00;
            12'b10110_0011101: DATA = 8'h00;
            12'b10110_0011110: DATA = 8'h00;
            12'b10110_0011111: DATA = 8'h00;
            12'b10110_0100000: DATA = 8'h00;
            12'b10110_0100001: DATA = 8'h00;
            12'b10110_0100010: DATA = 8'h00;
            12'b10110_0100011: DATA = 8'h00;
            12'b10110_0100100: DATA = 8'h00;
            12'b10110_0100101: DATA = 8'h00;
            12'b10110_0100110: DATA = 8'h00;
            12'b10110_0100111: DATA = 8'h00;
            12'b10110_0101000: DATA = 8'h00;
            12'b10110_0101001: DATA = 8'h00;
            12'b10110_0101010: DATA = 8'h00;
            12'b10110_0101011: DATA = 8'h00;
            12'b10110_0101100: DATA = 8'h00;
            12'b10110_0101101: DATA = 8'h00;
            12'b10110_0101110: DATA = 8'h00;
            12'b10110_0101111: DATA = 8'h00;
            12'b10110_0110000: DATA = 8'h00;
            12'b10110_0110001: DATA = 8'h00;
            12'b10110_0110010: DATA = 8'h00;
            12'b10110_0110011: DATA = 8'h00;
            12'b10110_0110100: DATA = 8'h00;
            12'b10110_0110101: DATA = 8'h00;
            12'b10110_0110110: DATA = 8'h00;
            12'b10110_0110111: DATA = 8'h00;
            12'b10110_0111000: DATA = 8'h00;
            12'b10110_0111001: DATA = 8'h00;
            12'b10110_0111010: DATA = 8'h00;
            12'b10110_0111011: DATA = 8'h00;
            12'b10110_0111100: DATA = 8'h00;
            12'b10110_0111101: DATA = 8'h00;
            12'b10110_0111110: DATA = 8'h00;
            12'b10110_0111111: DATA = 8'h00;
            12'b10110_1000000: DATA = 8'h00;
            12'b10110_1000001: DATA = 8'h00;
            12'b10110_1000010: DATA = 8'h00;
            12'b10110_1000011: DATA = 8'h00;
            12'b10110_1000100: DATA = 8'h00;
            12'b10110_1000101: DATA = 8'h00;
            12'b10110_1000110: DATA = 8'h00;
            12'b10110_1000111: DATA = 8'h00;
            12'b10110_1001000: DATA = 8'h00;
            12'b10110_1001001: DATA = 8'h00;
            12'b10110_1001010: DATA = 8'h00;
            12'b10110_1001011: DATA = 8'h00;
            12'b10110_1001100: DATA = 8'h00;
            12'b10110_1001101: DATA = 8'h00;
            12'b10110_1001110: DATA = 8'h00;
            12'b10110_1001111: DATA = 8'h00;
            // Row 23
            12'b10111_0000000: DATA = 8'h53;
            12'b10111_0000001: DATA = 8'h55;
            12'b10111_0000010: DATA = 8'h50;
            12'b10111_0000011: DATA = 8'h45;
            12'b10111_0000100: DATA = 8'h52;
            12'b10111_0000101: DATA = 8'h50;
            12'b10111_0000110: DATA = 8'h4F;
            12'b10111_0000111: DATA = 8'h53;
            12'b10111_0001000: DATA = 8'h49;
            12'b10111_0001001: DATA = 8'h54;
            12'b10111_0001010: DATA = 8'h49;
            12'b10111_0001011: DATA = 8'h4F;
            12'b10111_0001100: DATA = 8'h4E;
            12'b10111_0001101: DATA = 8'h00;
            12'b10111_0001110: DATA = 8'h4F;
            12'b10111_0001111: DATA = (SUPERPOSE == 1) ? 8'h4E : 8'h46;
            12'b10111_0010000: DATA = (SUPERPOSE == 1) ? 8'h00 : 8'h46;
            12'b10111_0010001: DATA = 8'h00;
            12'b10111_0010010: DATA = 8'h00;
            12'b10111_0010011: DATA = 8'h00;
            12'b10111_0010100: DATA = 8'h00;
            12'b10111_0010101: DATA = 8'h00;
            12'b10111_0010110: DATA = 8'h00;
            12'b10111_0010111: DATA = 8'h00;
            12'b10111_0011000: DATA = 8'h00;
            12'b10111_0011001: DATA = 8'h00;
            12'b10111_0011010: DATA = 8'h00;
            12'b10111_0011011: DATA = 8'h00;
            12'b10111_0011100: DATA = 8'h00;
            12'b10111_0011101: DATA = 8'h00;
            12'b10111_0011110: DATA = 8'h00;
            12'b10111_0011111: DATA = 8'h00;
            12'b10111_0100000: DATA = 8'h00;
            12'b10111_0100001: DATA = 8'h00;
            12'b10111_0100010: DATA = 8'h00;
            12'b10111_0100011: DATA = 8'h00;
            12'b10111_0100100: DATA = 8'h00;
            12'b10111_0100101: DATA = 8'h00;
            12'b10111_0100110: DATA = 8'h00;
            12'b10111_0100111: DATA = 8'h00;
            12'b10111_0101000: DATA = 8'h00;
            12'b10111_0101001: DATA = 8'h00;
            12'b10111_0101010: DATA = 8'h00;
            12'b10111_0101011: DATA = 8'h00;
            12'b10111_0101100: DATA = 8'h00;
            12'b10111_0101101: DATA = 8'h00;
            12'b10111_0101110: DATA = 8'h00;
            12'b10111_0101111: DATA = 8'h00;
            12'b10111_0110000: DATA = 8'h00;
            12'b10111_0110001: DATA = 8'h00;
            12'b10111_0110010: DATA = 8'h00;
            12'b10111_0110011: DATA = 8'h00;
            12'b10111_0110100: DATA = 8'h00;
            12'b10111_0110101: DATA = 8'h00;
            12'b10111_0110110: DATA = 8'h00;
            12'b10111_0110111: DATA = 8'h00;
            12'b10111_0111000: DATA = 8'h00;
            12'b10111_0111001: DATA = 8'h00;
            12'b10111_0111010: DATA = 8'h00;
            12'b10111_0111011: DATA = 8'h00;
            12'b10111_0111100: DATA = 8'h00;
            12'b10111_0111101: DATA = 8'h00;
            12'b10111_0111110: DATA = 8'h00;
            12'b10111_0111111: DATA = 8'h00;
            12'b10111_1000000: DATA = 8'h00;
            12'b10111_1000001: DATA = 8'h00;
            12'b10111_1000010: DATA = 8'h00;
            12'b10111_1000011: DATA = 8'h00;
            12'b10111_1000100: DATA = 8'h00;
            12'b10111_1000101: DATA = 8'h00;
            12'b10111_1000110: DATA = 8'h00;
            12'b10111_1000111: DATA = 8'h00;
            12'b10111_1001000: DATA = 8'h00;
            12'b10111_1001001: DATA = 8'h00;
            12'b10111_1001010: DATA = 8'h00;
            12'b10111_1001011: DATA = 8'h00;
            12'b10111_1001100: DATA = 8'h00;
            12'b10111_1001101: DATA = 8'h00;
            12'b10111_1001110: DATA = 8'h00;
            12'b10111_1001111: DATA = 8'h00;
            // Row 24
            12'b11000_0000000: DATA = 8'h00;
            12'b11000_0000001: DATA = 8'h00;
            12'b11000_0000010: DATA = 8'h00;
            12'b11000_0000011: DATA = 8'h00;
            12'b11000_0000100: DATA = 8'h00;
            12'b11000_0000101: DATA = 8'h00;
            12'b11000_0000110: DATA = 8'h00;
            12'b11000_0000111: DATA = 8'h00;
            12'b11000_0001000: DATA = 8'h00;
            12'b11000_0001001: DATA = 8'h00;
            12'b11000_0001010: DATA = 8'h00;
            12'b11000_0001011: DATA = 8'h00;
            12'b11000_0001100: DATA = 8'h00;
            12'b11000_0001101: DATA = 8'h00;
            12'b11000_0001110: DATA = 8'h00;
            12'b11000_0001111: DATA = 8'h00;
            12'b11000_0010000: DATA = 8'h00;
            12'b11000_0010001: DATA = 8'h00;
            12'b11000_0010010: DATA = 8'h00;
            12'b11000_0010011: DATA = 8'h00;
            12'b11000_0010100: DATA = 8'h00;
            12'b11000_0010101: DATA = 8'h00;
            12'b11000_0010110: DATA = 8'h00;
            12'b11000_0010111: DATA = 8'h00;
            12'b11000_0011000: DATA = 8'h00;
            12'b11000_0011001: DATA = 8'h00;
            12'b11000_0011010: DATA = 8'h00;
            12'b11000_0011011: DATA = 8'h00;
            12'b11000_0011100: DATA = 8'h00;
            12'b11000_0011101: DATA = 8'h00;
            12'b11000_0011110: DATA = 8'h00;
            12'b11000_0011111: DATA = 8'h00;
            12'b11000_0100000: DATA = 8'h00;
            12'b11000_0100001: DATA = 8'h00;
            12'b11000_0100010: DATA = 8'h00;
            12'b11000_0100011: DATA = 8'h00;
            12'b11000_0100100: DATA = 8'h00;
            12'b11000_0100101: DATA = 8'h00;
            12'b11000_0100110: DATA = 8'h00;
            12'b11000_0100111: DATA = 8'h00;
            12'b11000_0101000: DATA = 8'h00;
            12'b11000_0101001: DATA = 8'h00;
            12'b11000_0101010: DATA = 8'h00;
            12'b11000_0101011: DATA = 8'h00;
            12'b11000_0101100: DATA = 8'h00;
            12'b11000_0101101: DATA = 8'h00;
            12'b11000_0101110: DATA = 8'h00;
            12'b11000_0101111: DATA = 8'h00;
            12'b11000_0110000: DATA = 8'h00;
            12'b11000_0110001: DATA = 8'h00;
            12'b11000_0110010: DATA = 8'h00;
            12'b11000_0110011: DATA = 8'h00;
            12'b11000_0110100: DATA = 8'h00;
            12'b11000_0110101: DATA = 8'h00;
            12'b11000_0110110: DATA = 8'h00;
            12'b11000_0110111: DATA = 8'h00;
            12'b11000_0111000: DATA = 8'h00;
            12'b11000_0111001: DATA = 8'h00;
            12'b11000_0111010: DATA = 8'h00;
            12'b11000_0111011: DATA = 8'h00;
            12'b11000_0111100: DATA = 8'h00;
            12'b11000_0111101: DATA = 8'h00;
            12'b11000_0111110: DATA = 8'h00;
            12'b11000_0111111: DATA = 8'h00;
            12'b11000_1000000: DATA = 8'h00;
            12'b11000_1000001: DATA = 8'h00;
            12'b11000_1000010: DATA = 8'h00;
            12'b11000_1000011: DATA = 8'h00;
            12'b11000_1000100: DATA = 8'h00;
            12'b11000_1000101: DATA = 8'h00;
            12'b11000_1000110: DATA = 8'h00;
            12'b11000_1000111: DATA = 8'h00;
            12'b11000_1001000: DATA = 8'h00;
            12'b11000_1001001: DATA = 8'h00;
            12'b11000_1001010: DATA = 8'h00;
            12'b11000_1001011: DATA = 8'h00;
            12'b11000_1001100: DATA = 8'h00;
            12'b11000_1001101: DATA = 8'h00;
            12'b11000_1001110: DATA = 8'h00;
            12'b11000_1001111: DATA = 8'h00;
            // Row 25
            12'b11001_0000000: DATA = 8'h00;
            12'b11001_0000001: DATA = 8'h00;
            12'b11001_0000010: DATA = 8'h00;
            12'b11001_0000011: DATA = 8'h00;
            12'b11001_0000100: DATA = 8'h00;
            12'b11001_0000101: DATA = 8'h00;
            12'b11001_0000110: DATA = 8'h00;
            12'b11001_0000111: DATA = 8'h00;
            12'b11001_0001000: DATA = 8'h00;
            12'b11001_0001001: DATA = 8'h00;
            12'b11001_0001010: DATA = 8'h00;
            12'b11001_0001011: DATA = 8'h00;
            12'b11001_0001100: DATA = 8'h00;
            12'b11001_0001101: DATA = 8'h00;
            12'b11001_0001110: DATA = 8'h00;
            12'b11001_0001111: DATA = 8'h00;
            12'b11001_0010000: DATA = 8'h00;
            12'b11001_0010001: DATA = 8'h00;
            12'b11001_0010010: DATA = 8'h00;
            12'b11001_0010011: DATA = 8'h00;
            12'b11001_0010100: DATA = 8'h00;
            12'b11001_0010101: DATA = 8'h00;
            12'b11001_0010110: DATA = 8'h00;
            12'b11001_0010111: DATA = 8'h00;
            12'b11001_0011000: DATA = 8'h00;
            12'b11001_0011001: DATA = 8'h00;
            12'b11001_0011010: DATA = 8'h00;
            12'b11001_0011011: DATA = 8'h00;
            12'b11001_0011100: DATA = 8'h00;
            12'b11001_0011101: DATA = 8'h00;
            12'b11001_0011110: DATA = 8'h00;
            12'b11001_0011111: DATA = 8'h00;
            12'b11001_0100000: DATA = 8'h00;
            12'b11001_0100001: DATA = 8'h00;
            12'b11001_0100010: DATA = 8'h00;
            12'b11001_0100011: DATA = 8'h00;
            12'b11001_0100100: DATA = 8'h00;
            12'b11001_0100101: DATA = 8'h00;
            12'b11001_0100110: DATA = 8'h00;
            12'b11001_0100111: DATA = 8'h00;
            12'b11001_0101000: DATA = 8'h00;
            12'b11001_0101001: DATA = 8'h00;
            12'b11001_0101010: DATA = 8'h00;
            12'b11001_0101011: DATA = 8'h00;
            12'b11001_0101100: DATA = 8'h00;
            12'b11001_0101101: DATA = 8'h00;
            12'b11001_0101110: DATA = 8'h00;
            12'b11001_0101111: DATA = 8'h00;
            12'b11001_0110000: DATA = 8'h00;
            12'b11001_0110001: DATA = 8'h00;
            12'b11001_0110010: DATA = 8'h00;
            12'b11001_0110011: DATA = 8'h00;
            12'b11001_0110100: DATA = 8'h00;
            12'b11001_0110101: DATA = 8'h00;
            12'b11001_0110110: DATA = 8'h00;
            12'b11001_0110111: DATA = 8'h00;
            12'b11001_0111000: DATA = 8'h00;
            12'b11001_0111001: DATA = 8'h00;
            12'b11001_0111010: DATA = 8'h00;
            12'b11001_0111011: DATA = 8'h00;
            12'b11001_0111100: DATA = 8'h00;
            12'b11001_0111101: DATA = 8'h00;
            12'b11001_0111110: DATA = 8'h00;
            12'b11001_0111111: DATA = 8'h00;
            12'b11001_1000000: DATA = 8'h00;
            12'b11001_1000001: DATA = 8'h00;
            12'b11001_1000010: DATA = 8'h00;
            12'b11001_1000011: DATA = 8'h00;
            12'b11001_1000100: DATA = 8'h00;
            12'b11001_1000101: DATA = 8'h00;
            12'b11001_1000110: DATA = 8'h00;
            12'b11001_1000111: DATA = 8'h00;
            12'b11001_1001000: DATA = 8'h00;
            12'b11001_1001001: DATA = 8'h00;
            12'b11001_1001010: DATA = 8'h00;
            12'b11001_1001011: DATA = 8'h00;
            12'b11001_1001100: DATA = 8'h00;
            12'b11001_1001101: DATA = 8'h00;
            12'b11001_1001110: DATA = 8'h00;
            12'b11001_1001111: DATA = 8'h00;
            // Row 26
            12'b11010_0000000: DATA = 8'h00;
            12'b11010_0000001: DATA = 8'h00;
            12'b11010_0000010: DATA = 8'h00;
            12'b11010_0000011: DATA = 8'h00;
            12'b11010_0000100: DATA = 8'h00;
            12'b11010_0000101: DATA = 8'h00;
            12'b11010_0000110: DATA = 8'h00;
            12'b11010_0000111: DATA = 8'h00;
            12'b11010_0001000: DATA = 8'h00;
            12'b11010_0001001: DATA = 8'h00;
            12'b11010_0001010: DATA = 8'h00;
            12'b11010_0001011: DATA = 8'h00;
            12'b11010_0001100: DATA = 8'h00;
            12'b11010_0001101: DATA = 8'h00;
            12'b11010_0001110: DATA = 8'h00;
            12'b11010_0001111: DATA = 8'h00;
            12'b11010_0010000: DATA = 8'h00;
            12'b11010_0010001: DATA = 8'h00;
            12'b11010_0010010: DATA = 8'h00;
            12'b11010_0010011: DATA = 8'h00;
            12'b11010_0010100: DATA = 8'h00;
            12'b11010_0010101: DATA = 8'h00;
            12'b11010_0010110: DATA = 8'h00;
            12'b11010_0010111: DATA = 8'h00;
            12'b11010_0011000: DATA = 8'h00;
            12'b11010_0011001: DATA = 8'h00;
            12'b11010_0011010: DATA = 8'h00;
            12'b11010_0011011: DATA = 8'h00;
            12'b11010_0011100: DATA = 8'h00;
            12'b11010_0011101: DATA = 8'h00;
            12'b11010_0011110: DATA = 8'h00;
            12'b11010_0011111: DATA = 8'h00;
            12'b11010_0100000: DATA = 8'h00;
            12'b11010_0100001: DATA = 8'h00;
            12'b11010_0100010: DATA = 8'h00;
            12'b11010_0100011: DATA = 8'h00;
            12'b11010_0100100: DATA = 8'h00;
            12'b11010_0100101: DATA = 8'h00;
            12'b11010_0100110: DATA = 8'h00;
            12'b11010_0100111: DATA = 8'h00;
            12'b11010_0101000: DATA = 8'h00;
            12'b11010_0101001: DATA = 8'h00;
            12'b11010_0101010: DATA = 8'h00;
            12'b11010_0101011: DATA = 8'h00;
            12'b11010_0101100: DATA = 8'h00;
            12'b11010_0101101: DATA = 8'h00;
            12'b11010_0101110: DATA = 8'h00;
            12'b11010_0101111: DATA = 8'h00;
            12'b11010_0110000: DATA = 8'h00;
            12'b11010_0110001: DATA = 8'h00;
            12'b11010_0110010: DATA = 8'h00;
            12'b11010_0110011: DATA = 8'h00;
            12'b11010_0110100: DATA = 8'h00;
            12'b11010_0110101: DATA = 8'h00;
            12'b11010_0110110: DATA = 8'h00;
            12'b11010_0110111: DATA = 8'h00;
            12'b11010_0111000: DATA = 8'h00;
            12'b11010_0111001: DATA = 8'h00;
            12'b11010_0111010: DATA = 8'h00;
            12'b11010_0111011: DATA = 8'h00;
            12'b11010_0111100: DATA = 8'h00;
            12'b11010_0111101: DATA = 8'h00;
            12'b11010_0111110: DATA = 8'h00;
            12'b11010_0111111: DATA = 8'h00;
            12'b11010_1000000: DATA = 8'h00;
            12'b11010_1000001: DATA = 8'h00;
            12'b11010_1000010: DATA = 8'h00;
            12'b11010_1000011: DATA = 8'h00;
            12'b11010_1000100: DATA = 8'h00;
            12'b11010_1000101: DATA = 8'h00;
            12'b11010_1000110: DATA = 8'h00;
            12'b11010_1000111: DATA = 8'h00;
            12'b11010_1001000: DATA = 8'h00;
            12'b11010_1001001: DATA = 8'h00;
            12'b11010_1001010: DATA = 8'h00;
            12'b11010_1001011: DATA = 8'h00;
            12'b11010_1001100: DATA = 8'h00;
            12'b11010_1001101: DATA = 8'h00;
            12'b11010_1001110: DATA = 8'h00;
            12'b11010_1001111: DATA = 8'h00;
            // Row 27
            12'b11011_0000000: DATA = 8'h00;
            12'b11011_0000001: DATA = 8'h00;
            12'b11011_0000010: DATA = 8'h00;
            12'b11011_0000011: DATA = 8'h00;
            12'b11011_0000100: DATA = 8'h00;
            12'b11011_0000101: DATA = 8'h00;
            12'b11011_0000110: DATA = 8'h00;
            12'b11011_0000111: DATA = 8'h00;
            12'b11011_0001000: DATA = 8'h00;
            12'b11011_0001001: DATA = 8'h00;
            12'b11011_0001010: DATA = 8'h00;
            12'b11011_0001011: DATA = 8'h00;
            12'b11011_0001100: DATA = 8'h00;
            12'b11011_0001101: DATA = 8'h00;
            12'b11011_0001110: DATA = 8'h00;
            12'b11011_0001111: DATA = 8'h00;
            12'b11011_0010000: DATA = 8'h00;
            12'b11011_0010001: DATA = 8'h00;
            12'b11011_0010010: DATA = 8'h00;
            12'b11011_0010011: DATA = 8'h00;
            12'b11011_0010100: DATA = 8'h00;
            12'b11011_0010101: DATA = 8'h00;
            12'b11011_0010110: DATA = 8'h00;
            12'b11011_0010111: DATA = 8'h00;
            12'b11011_0011000: DATA = 8'h00;
            12'b11011_0011001: DATA = 8'h00;
            12'b11011_0011010: DATA = 8'h00;
            12'b11011_0011011: DATA = 8'h00;
            12'b11011_0011100: DATA = 8'h00;
            12'b11011_0011101: DATA = 8'h00;
            12'b11011_0011110: DATA = 8'h00;
            12'b11011_0011111: DATA = 8'h00;
            12'b11011_0100000: DATA = 8'h00;
            12'b11011_0100001: DATA = 8'h00;
            12'b11011_0100010: DATA = 8'h00;
            12'b11011_0100011: DATA = 8'h00;
            12'b11011_0100100: DATA = 8'h00;
            12'b11011_0100101: DATA = 8'h00;
            12'b11011_0100110: DATA = 8'h00;
            12'b11011_0100111: DATA = 8'h00;
            12'b11011_0101000: DATA = 8'h00;
            12'b11011_0101001: DATA = 8'h00;
            12'b11011_0101010: DATA = 8'h00;
            12'b11011_0101011: DATA = 8'h00;
            12'b11011_0101100: DATA = 8'h00;
            12'b11011_0101101: DATA = 8'h00;
            12'b11011_0101110: DATA = 8'h00;
            12'b11011_0101111: DATA = 8'h00;
            12'b11011_0110000: DATA = 8'h00;
            12'b11011_0110001: DATA = 8'h00;
            12'b11011_0110010: DATA = 8'h00;
            12'b11011_0110011: DATA = 8'h00;
            12'b11011_0110100: DATA = 8'h00;
            12'b11011_0110101: DATA = 8'h00;
            12'b11011_0110110: DATA = 8'h00;
            12'b11011_0110111: DATA = 8'h00;
            12'b11011_0111000: DATA = 8'h00;
            12'b11011_0111001: DATA = 8'h00;
            12'b11011_0111010: DATA = 8'h00;
            12'b11011_0111011: DATA = 8'h00;
            12'b11011_0111100: DATA = 8'h00;
            12'b11011_0111101: DATA = 8'h00;
            12'b11011_0111110: DATA = 8'h00;
            12'b11011_0111111: DATA = 8'h00;
            12'b11011_1000000: DATA = 8'h00;
            12'b11011_1000001: DATA = 8'h00;
            12'b11011_1000010: DATA = 8'h00;
            12'b11011_1000011: DATA = 8'h00;
            12'b11011_1000100: DATA = 8'h00;
            12'b11011_1000101: DATA = 8'h00;
            12'b11011_1000110: DATA = 8'h00;
            12'b11011_1000111: DATA = 8'h00;
            12'b11011_1001000: DATA = 8'h00;
            12'b11011_1001001: DATA = 8'h00;
            12'b11011_1001010: DATA = 8'h00;
            12'b11011_1001011: DATA = 8'h00;
            12'b11011_1001100: DATA = 8'h00;
            12'b11011_1001101: DATA = 8'h00;
            12'b11011_1001110: DATA = 8'h00;
            12'b11011_1001111: DATA = 8'h00;
            // Row 28
            12'b11100_0000000: DATA = 8'h00;
            12'b11100_0000001: DATA = 8'h00;
            12'b11100_0000010: DATA = 8'h00;
            12'b11100_0000011: DATA = 8'h00;
            12'b11100_0000100: DATA = 8'h00;
            12'b11100_0000101: DATA = 8'h00;
            12'b11100_0000110: DATA = 8'h00;
            12'b11100_0000111: DATA = 8'h00;
            12'b11100_0001000: DATA = 8'h00;
            12'b11100_0001001: DATA = 8'h00;
            12'b11100_0001010: DATA = 8'h00;
            12'b11100_0001011: DATA = 8'h00;
            12'b11100_0001100: DATA = 8'h00;
            12'b11100_0001101: DATA = 8'h00;
            12'b11100_0001110: DATA = 8'h00;
            12'b11100_0001111: DATA = 8'h00;
            12'b11100_0010000: DATA = 8'h00;
            12'b11100_0010001: DATA = 8'h00;
            12'b11100_0010010: DATA = 8'h00;
            12'b11100_0010011: DATA = 8'h00;
            12'b11100_0010100: DATA = 8'h00;
            12'b11100_0010101: DATA = 8'h00;
            12'b11100_0010110: DATA = 8'h00;
            12'b11100_0010111: DATA = 8'h00;
            12'b11100_0011000: DATA = 8'h00;
            12'b11100_0011001: DATA = 8'h00;
            12'b11100_0011010: DATA = 8'h00;
            12'b11100_0011011: DATA = 8'h00;
            12'b11100_0011100: DATA = 8'h00;
            12'b11100_0011101: DATA = 8'h00;
            12'b11100_0011110: DATA = 8'h00;
            12'b11100_0011111: DATA = 8'h00;
            12'b11100_0100000: DATA = 8'h00;
            12'b11100_0100001: DATA = 8'h00;
            12'b11100_0100010: DATA = 8'h00;
            12'b11100_0100011: DATA = 8'h00;
            12'b11100_0100100: DATA = 8'h00;
            12'b11100_0100101: DATA = 8'h00;
            12'b11100_0100110: DATA = 8'h00;
            12'b11100_0100111: DATA = 8'h00;
            12'b11100_0101000: DATA = 8'h00;
            12'b11100_0101001: DATA = 8'h00;
            12'b11100_0101010: DATA = 8'h00;
            12'b11100_0101011: DATA = 8'h00;
            12'b11100_0101100: DATA = 8'h00;
            12'b11100_0101101: DATA = 8'h00;
            12'b11100_0101110: DATA = 8'h00;
            12'b11100_0101111: DATA = 8'h00;
            12'b11100_0110000: DATA = 8'h00;
            12'b11100_0110001: DATA = 8'h00;
            12'b11100_0110010: DATA = 8'h00;
            12'b11100_0110011: DATA = 8'h00;
            12'b11100_0110100: DATA = 8'h00;
            12'b11100_0110101: DATA = 8'h00;
            12'b11100_0110110: DATA = 8'h00;
            12'b11100_0110111: DATA = 8'h00;
            12'b11100_0111000: DATA = 8'h00;
            12'b11100_0111001: DATA = 8'h00;
            12'b11100_0111010: DATA = 8'h00;
            12'b11100_0111011: DATA = 8'h00;
            12'b11100_0111100: DATA = 8'h00;
            12'b11100_0111101: DATA = 8'h00;
            12'b11100_0111110: DATA = 8'h00;
            12'b11100_0111111: DATA = 8'h00;
            12'b11100_1000000: DATA = 8'h00;
            12'b11100_1000001: DATA = 8'h00;
            12'b11100_1000010: DATA = 8'h00;
            12'b11100_1000011: DATA = 8'h00;
            12'b11100_1000100: DATA = 8'h00;
            12'b11100_1000101: DATA = 8'h00;
            12'b11100_1000110: DATA = 8'h00;
            12'b11100_1000111: DATA = 8'h00;
            12'b11100_1001000: DATA = 8'h00;
            12'b11100_1001001: DATA = 8'h00;
            12'b11100_1001010: DATA = 8'h00;
            12'b11100_1001011: DATA = 8'h00;
            12'b11100_1001100: DATA = 8'h00;
            12'b11100_1001101: DATA = 8'h00;
            12'b11100_1001110: DATA = 8'h00;
            12'b11100_1001111: DATA = 8'h00;
            // Row 29
            12'b11101_0000000: DATA = 8'h00;
            12'b11101_0000001: DATA = 8'h00;
            12'b11101_0000010: DATA = 8'h00;
            12'b11101_0000011: DATA = 8'h00;
            12'b11101_0000100: DATA = 8'h00;
            12'b11101_0000101: DATA = 8'h00;
            12'b11101_0000110: DATA = 8'h00;
            12'b11101_0000111: DATA = 8'h00;
            12'b11101_0001000: DATA = 8'h00;
            12'b11101_0001001: DATA = 8'h00;
            12'b11101_0001010: DATA = 8'h00;
            12'b11101_0001011: DATA = 8'h00;
            12'b11101_0001100: DATA = 8'h00;
            12'b11101_0001101: DATA = 8'h00;
            12'b11101_0001110: DATA = 8'h00;
            12'b11101_0001111: DATA = 8'h00;
            12'b11101_0010000: DATA = 8'h00;
            12'b11101_0010001: DATA = 8'h00;
            12'b11101_0010010: DATA = 8'h00;
            12'b11101_0010011: DATA = 8'h00;
            12'b11101_0010100: DATA = 8'h00;
            12'b11101_0010101: DATA = 8'h00;
            12'b11101_0010110: DATA = 8'h00;
            12'b11101_0010111: DATA = 8'h00;
            12'b11101_0011000: DATA = 8'h00;
            12'b11101_0011001: DATA = 8'h00;
            12'b11101_0011010: DATA = 8'h00;
            12'b11101_0011011: DATA = 8'h00;
            12'b11101_0011100: DATA = 8'h00;
            12'b11101_0011101: DATA = 8'h00;
            12'b11101_0011110: DATA = 8'h00;
            12'b11101_0011111: DATA = 8'h00;
            12'b11101_0100000: DATA = 8'h00;
            12'b11101_0100001: DATA = 8'h00;
            12'b11101_0100010: DATA = 8'h00;
            12'b11101_0100011: DATA = 8'h00;
            12'b11101_0100100: DATA = 8'h00;
            12'b11101_0100101: DATA = 8'h00;
            12'b11101_0100110: DATA = 8'h00;
            12'b11101_0100111: DATA = 8'h00;
            12'b11101_0101000: DATA = 8'h00;
            12'b11101_0101001: DATA = 8'h00;
            12'b11101_0101010: DATA = 8'h00;
            12'b11101_0101011: DATA = 8'h00;
            12'b11101_0101100: DATA = 8'h00;
            12'b11101_0101101: DATA = 8'h00;
            12'b11101_0101110: DATA = 8'h00;
            12'b11101_0101111: DATA = 8'h00;
            12'b11101_0110000: DATA = 8'h00;
            12'b11101_0110001: DATA = 8'h00;
            12'b11101_0110010: DATA = 8'h00;
            12'b11101_0110011: DATA = 8'h00;
            12'b11101_0110100: DATA = 8'h00;
            12'b11101_0110101: DATA = 8'h00;
            12'b11101_0110110: DATA = 8'h00;
            12'b11101_0110111: DATA = 8'h00;
            12'b11101_0111000: DATA = 8'h00;
            12'b11101_0111001: DATA = 8'h00;
            12'b11101_0111010: DATA = 8'h00;
            12'b11101_0111011: DATA = 8'h00;
            12'b11101_0111100: DATA = 8'h00;
            12'b11101_0111101: DATA = 8'h00;
            12'b11101_0111110: DATA = 8'h00;
            12'b11101_0111111: DATA = 8'h00;
            12'b11101_1000000: DATA = 8'h00;
            12'b11101_1000001: DATA = 8'h00;
            12'b11101_1000010: DATA = 8'h00;
            12'b11101_1000011: DATA = 8'h00;
            12'b11101_1000100: DATA = 8'h00;
            12'b11101_1000101: DATA = 8'h00;
            12'b11101_1000110: DATA = 8'h00;
            12'b11101_1000111: DATA = 8'h00;
            12'b11101_1001000: DATA = 8'h00;
            12'b11101_1001001: DATA = 8'h00;
            12'b11101_1001010: DATA = 8'h00;
            12'b11101_1001011: DATA = 8'h00;
            12'b11101_1001100: DATA = 8'h00;
            12'b11101_1001101: DATA = 8'h00;
            12'b11101_1001110: DATA = 8'h00;
            12'b11101_1001111: DATA = 8'h00;
            default: DATA = 8'h00;
        endcase
    end
endmodule
