`timescale 1ns / 1ps

module display_rom(
    input CLK,
    input [7:0] CHAR,
    input [3:0] ROW,
    input [2:0] COL,
    output reg DATA
    );
    
    reg [7:0] CHAR_REG;
    reg [3:0] ROW_REG;
    reg [2:0] COL_REG;
    
    always @ (posedge CLK) begin
        CHAR_REG <= CHAR;
        ROW_REG <= ROW;
        COL_REG <= COL;
    end
    
    always @ (*) begin
        case ({CHAR_REG, ROW_REG, COL_REG})
            // ' Row 0
            15'b00100111_0000_000: DATA = 1'b0;
            15'b00100111_0000_001: DATA = 1'b0;
            15'b00100111_0000_010: DATA = 1'b0;
            15'b00100111_0000_011: DATA = 1'b0;
            15'b00100111_0000_100: DATA = 1'b0;
            15'b00100111_0000_101: DATA = 1'b0;
            15'b00100111_0000_110: DATA = 1'b0;
            15'b00100111_0000_111: DATA = 1'b0;
            // ' Row 1
            15'b00100111_0001_000: DATA = 1'b0;
            15'b00100111_0001_001: DATA = 1'b0;
            15'b00100111_0001_010: DATA = 1'b0;
            15'b00100111_0001_011: DATA = 1'b0;
            15'b00100111_0001_100: DATA = 1'b0;
            15'b00100111_0001_101: DATA = 1'b0;
            15'b00100111_0001_110: DATA = 1'b0;
            15'b00100111_0001_111: DATA = 1'b0;
            // ' Row 2
            15'b00100111_0010_000: DATA = 1'b0;
            15'b00100111_0010_001: DATA = 1'b0;
            15'b00100111_0010_010: DATA = 1'b0;
            15'b00100111_0010_011: DATA = 1'b0;
            15'b00100111_0010_100: DATA = 1'b0;
            15'b00100111_0010_101: DATA = 1'b0;
            15'b00100111_0010_110: DATA = 1'b0;
            15'b00100111_0010_111: DATA = 1'b0;
            // ' Row 3
            15'b00100111_0011_000: DATA = 1'b0;
            15'b00100111_0011_001: DATA = 1'b0;
            15'b00100111_0011_010: DATA = 1'b1;
            15'b00100111_0011_011: DATA = 1'b1;
            15'b00100111_0011_100: DATA = 1'b0;
            15'b00100111_0011_101: DATA = 1'b0;
            15'b00100111_0011_110: DATA = 1'b0;
            15'b00100111_0011_111: DATA = 1'b0;
            // ' Row 4
            15'b00100111_0100_000: DATA = 1'b0;
            15'b00100111_0100_001: DATA = 1'b0;
            15'b00100111_0100_010: DATA = 1'b1;
            15'b00100111_0100_011: DATA = 1'b1;
            15'b00100111_0100_100: DATA = 1'b0;
            15'b00100111_0100_101: DATA = 1'b0;
            15'b00100111_0100_110: DATA = 1'b0;
            15'b00100111_0100_111: DATA = 1'b0;
            // ' Row 5
            15'b00100111_0101_000: DATA = 1'b0;
            15'b00100111_0101_001: DATA = 1'b1;
            15'b00100111_0101_010: DATA = 1'b1;
            15'b00100111_0101_011: DATA = 1'b0;
            15'b00100111_0101_100: DATA = 1'b0;
            15'b00100111_0101_101: DATA = 1'b0;
            15'b00100111_0101_110: DATA = 1'b0;
            15'b00100111_0101_111: DATA = 1'b0;
            // ' Row 6
            15'b00100111_0110_000: DATA = 1'b0;
            15'b00100111_0110_001: DATA = 1'b0;
            15'b00100111_0110_010: DATA = 1'b0;
            15'b00100111_0110_011: DATA = 1'b0;
            15'b00100111_0110_100: DATA = 1'b0;
            15'b00100111_0110_101: DATA = 1'b0;
            15'b00100111_0110_110: DATA = 1'b0;
            15'b00100111_0110_111: DATA = 1'b0;
            // ' Row 7
            15'b00100111_0111_000: DATA = 1'b0;
            15'b00100111_0111_001: DATA = 1'b0;
            15'b00100111_0111_010: DATA = 1'b0;
            15'b00100111_0111_011: DATA = 1'b0;
            15'b00100111_0111_100: DATA = 1'b0;
            15'b00100111_0111_101: DATA = 1'b0;
            15'b00100111_0111_110: DATA = 1'b0;
            15'b00100111_0111_111: DATA = 1'b0;
            // ' Row 8
            15'b00100111_1000_000: DATA = 1'b0;
            15'b00100111_1000_001: DATA = 1'b0;
            15'b00100111_1000_010: DATA = 1'b0;
            15'b00100111_1000_011: DATA = 1'b0;
            15'b00100111_1000_100: DATA = 1'b0;
            15'b00100111_1000_101: DATA = 1'b0;
            15'b00100111_1000_110: DATA = 1'b0;
            15'b00100111_1000_111: DATA = 1'b0;
            // ' Row 9
            15'b00100111_1001_000: DATA = 1'b0;
            15'b00100111_1001_001: DATA = 1'b0;
            15'b00100111_1001_010: DATA = 1'b0;
            15'b00100111_1001_011: DATA = 1'b0;
            15'b00100111_1001_100: DATA = 1'b0;
            15'b00100111_1001_101: DATA = 1'b0;
            15'b00100111_1001_110: DATA = 1'b0;
            15'b00100111_1001_111: DATA = 1'b0;
            // ' Row 10
            15'b00100111_1010_000: DATA = 1'b0;
            15'b00100111_1010_001: DATA = 1'b0;
            15'b00100111_1010_010: DATA = 1'b0;
            15'b00100111_1010_011: DATA = 1'b0;
            15'b00100111_1010_100: DATA = 1'b0;
            15'b00100111_1010_101: DATA = 1'b0;
            15'b00100111_1010_110: DATA = 1'b0;
            15'b00100111_1010_111: DATA = 1'b0;
            // ' Row 11
            15'b00100111_1011_000: DATA = 1'b0;
            15'b00100111_1011_001: DATA = 1'b0;
            15'b00100111_1011_010: DATA = 1'b0;
            15'b00100111_1011_011: DATA = 1'b0;
            15'b00100111_1011_100: DATA = 1'b0;
            15'b00100111_1011_101: DATA = 1'b0;
            15'b00100111_1011_110: DATA = 1'b0;
            15'b00100111_1011_111: DATA = 1'b0;
            // ' Row 12
            15'b00100111_1100_000: DATA = 1'b0;
            15'b00100111_1100_001: DATA = 1'b0;
            15'b00100111_1100_010: DATA = 1'b0;
            15'b00100111_1100_011: DATA = 1'b0;
            15'b00100111_1100_100: DATA = 1'b0;
            15'b00100111_1100_101: DATA = 1'b0;
            15'b00100111_1100_110: DATA = 1'b0;
            15'b00100111_1100_111: DATA = 1'b0;
            // ' Row 13
            15'b00100111_1101_000: DATA = 1'b0;
            15'b00100111_1101_001: DATA = 1'b0;
            15'b00100111_1101_010: DATA = 1'b0;
            15'b00100111_1101_011: DATA = 1'b0;
            15'b00100111_1101_100: DATA = 1'b0;
            15'b00100111_1101_101: DATA = 1'b0;
            15'b00100111_1101_110: DATA = 1'b0;
            15'b00100111_1101_111: DATA = 1'b0;
            // ' Row 14
            15'b00100111_1110_000: DATA = 1'b0;
            15'b00100111_1110_001: DATA = 1'b0;
            15'b00100111_1110_010: DATA = 1'b0;
            15'b00100111_1110_011: DATA = 1'b0;
            15'b00100111_1110_100: DATA = 1'b0;
            15'b00100111_1110_101: DATA = 1'b0;
            15'b00100111_1110_110: DATA = 1'b0;
            15'b00100111_1110_111: DATA = 1'b0;
            // ' Row 15
            15'b00100111_1111_000: DATA = 1'b0;
            15'b00100111_1111_001: DATA = 1'b0;
            15'b00100111_1111_010: DATA = 1'b0;
            15'b00100111_1111_011: DATA = 1'b0;
            15'b00100111_1111_100: DATA = 1'b0;
            15'b00100111_1111_101: DATA = 1'b0;
            15'b00100111_1111_110: DATA = 1'b0;
            15'b00100111_1111_111: DATA = 1'b0;
            // - Row 0
            15'b00101101_0000_000: DATA = 1'b0;
            15'b00101101_0000_001: DATA = 1'b0;
            15'b00101101_0000_010: DATA = 1'b0;
            15'b00101101_0000_011: DATA = 1'b0;
            15'b00101101_0000_100: DATA = 1'b0;
            15'b00101101_0000_101: DATA = 1'b0;
            15'b00101101_0000_110: DATA = 1'b0;
            15'b00101101_0000_111: DATA = 1'b0;
            // - Row 1
            15'b00101101_0001_000: DATA = 1'b0;
            15'b00101101_0001_001: DATA = 1'b0;
            15'b00101101_0001_010: DATA = 1'b0;
            15'b00101101_0001_011: DATA = 1'b0;
            15'b00101101_0001_100: DATA = 1'b0;
            15'b00101101_0001_101: DATA = 1'b0;
            15'b00101101_0001_110: DATA = 1'b0;
            15'b00101101_0001_111: DATA = 1'b0;
            // - Row 2
            15'b00101101_0010_000: DATA = 1'b0;
            15'b00101101_0010_001: DATA = 1'b0;
            15'b00101101_0010_010: DATA = 1'b0;
            15'b00101101_0010_011: DATA = 1'b0;
            15'b00101101_0010_100: DATA = 1'b0;
            15'b00101101_0010_101: DATA = 1'b0;
            15'b00101101_0010_110: DATA = 1'b0;
            15'b00101101_0010_111: DATA = 1'b0;
            // - Row 3
            15'b00101101_0011_000: DATA = 1'b0;
            15'b00101101_0011_001: DATA = 1'b0;
            15'b00101101_0011_010: DATA = 1'b0;
            15'b00101101_0011_011: DATA = 1'b0;
            15'b00101101_0011_100: DATA = 1'b0;
            15'b00101101_0011_101: DATA = 1'b0;
            15'b00101101_0011_110: DATA = 1'b0;
            15'b00101101_0011_111: DATA = 1'b0;
            // - Row 4
            15'b00101101_0100_000: DATA = 1'b0;
            15'b00101101_0100_001: DATA = 1'b0;
            15'b00101101_0100_010: DATA = 1'b0;
            15'b00101101_0100_011: DATA = 1'b0;
            15'b00101101_0100_100: DATA = 1'b0;
            15'b00101101_0100_101: DATA = 1'b0;
            15'b00101101_0100_110: DATA = 1'b0;
            15'b00101101_0100_111: DATA = 1'b0;
            // - Row 5
            15'b00101101_0101_000: DATA = 1'b0;
            15'b00101101_0101_001: DATA = 1'b0;
            15'b00101101_0101_010: DATA = 1'b0;
            15'b00101101_0101_011: DATA = 1'b0;
            15'b00101101_0101_100: DATA = 1'b0;
            15'b00101101_0101_101: DATA = 1'b0;
            15'b00101101_0101_110: DATA = 1'b0;
            15'b00101101_0101_111: DATA = 1'b0;
            // - Row 6
            15'b00101101_0110_000: DATA = 1'b0;
            15'b00101101_0110_001: DATA = 1'b0;
            15'b00101101_0110_010: DATA = 1'b0;
            15'b00101101_0110_011: DATA = 1'b0;
            15'b00101101_0110_100: DATA = 1'b0;
            15'b00101101_0110_101: DATA = 1'b0;
            15'b00101101_0110_110: DATA = 1'b0;
            15'b00101101_0110_111: DATA = 1'b0;
            // - Row 7
            15'b00101101_0111_000: DATA = 1'b0;
            15'b00101101_0111_001: DATA = 1'b1;
            15'b00101101_0111_010: DATA = 1'b1;
            15'b00101101_0111_011: DATA = 1'b1;
            15'b00101101_0111_100: DATA = 1'b1;
            15'b00101101_0111_101: DATA = 1'b1;
            15'b00101101_0111_110: DATA = 1'b0;
            15'b00101101_0111_111: DATA = 1'b0;
            // - Row 8
            15'b00101101_1000_000: DATA = 1'b0;
            15'b00101101_1000_001: DATA = 1'b1;
            15'b00101101_1000_010: DATA = 1'b1;
            15'b00101101_1000_011: DATA = 1'b1;
            15'b00101101_1000_100: DATA = 1'b1;
            15'b00101101_1000_101: DATA = 1'b1;
            15'b00101101_1000_110: DATA = 1'b0;
            15'b00101101_1000_111: DATA = 1'b0;
            // - Row 9
            15'b00101101_1001_000: DATA = 1'b0;
            15'b00101101_1001_001: DATA = 1'b0;
            15'b00101101_1001_010: DATA = 1'b0;
            15'b00101101_1001_011: DATA = 1'b0;
            15'b00101101_1001_100: DATA = 1'b0;
            15'b00101101_1001_101: DATA = 1'b0;
            15'b00101101_1001_110: DATA = 1'b0;
            15'b00101101_1001_111: DATA = 1'b0;
            // - Row 10
            15'b00101101_1010_000: DATA = 1'b0;
            15'b00101101_1010_001: DATA = 1'b0;
            15'b00101101_1010_010: DATA = 1'b0;
            15'b00101101_1010_011: DATA = 1'b0;
            15'b00101101_1010_100: DATA = 1'b0;
            15'b00101101_1010_101: DATA = 1'b0;
            15'b00101101_1010_110: DATA = 1'b0;
            15'b00101101_1010_111: DATA = 1'b0;
            // - Row 11
            15'b00101101_1011_000: DATA = 1'b0;
            15'b00101101_1011_001: DATA = 1'b0;
            15'b00101101_1011_010: DATA = 1'b0;
            15'b00101101_1011_011: DATA = 1'b0;
            15'b00101101_1011_100: DATA = 1'b0;
            15'b00101101_1011_101: DATA = 1'b0;
            15'b00101101_1011_110: DATA = 1'b0;
            15'b00101101_1011_111: DATA = 1'b0;
            // - Row 12
            15'b00101101_1100_000: DATA = 1'b0;
            15'b00101101_1100_001: DATA = 1'b0;
            15'b00101101_1100_010: DATA = 1'b0;
            15'b00101101_1100_011: DATA = 1'b0;
            15'b00101101_1100_100: DATA = 1'b0;
            15'b00101101_1100_101: DATA = 1'b0;
            15'b00101101_1100_110: DATA = 1'b0;
            15'b00101101_1100_111: DATA = 1'b0;
            // - Row 13
            15'b00101101_1101_000: DATA = 1'b0;
            15'b00101101_1101_001: DATA = 1'b0;
            15'b00101101_1101_010: DATA = 1'b0;
            15'b00101101_1101_011: DATA = 1'b0;
            15'b00101101_1101_100: DATA = 1'b0;
            15'b00101101_1101_101: DATA = 1'b0;
            15'b00101101_1101_110: DATA = 1'b0;
            15'b00101101_1101_111: DATA = 1'b0;
            // - Row 14
            15'b00101101_1110_000: DATA = 1'b0;
            15'b00101101_1110_001: DATA = 1'b0;
            15'b00101101_1110_010: DATA = 1'b0;
            15'b00101101_1110_011: DATA = 1'b0;
            15'b00101101_1110_100: DATA = 1'b0;
            15'b00101101_1110_101: DATA = 1'b0;
            15'b00101101_1110_110: DATA = 1'b0;
            15'b00101101_1110_111: DATA = 1'b0;
            // - Row 15
            15'b00101101_1111_000: DATA = 1'b0;
            15'b00101101_1111_001: DATA = 1'b0;
            15'b00101101_1111_010: DATA = 1'b0;
            15'b00101101_1111_011: DATA = 1'b0;
            15'b00101101_1111_100: DATA = 1'b0;
            15'b00101101_1111_101: DATA = 1'b0;
            15'b00101101_1111_110: DATA = 1'b0;
            15'b00101101_1111_111: DATA = 1'b0;
            // . Row 0
            15'b00101110_0000_000: DATA = 1'b0;
            15'b00101110_0000_001: DATA = 1'b0;
            15'b00101110_0000_010: DATA = 1'b0;
            15'b00101110_0000_011: DATA = 1'b0;
            15'b00101110_0000_100: DATA = 1'b0;
            15'b00101110_0000_101: DATA = 1'b0;
            15'b00101110_0000_110: DATA = 1'b0;
            15'b00101110_0000_111: DATA = 1'b0;
            // . Row 1
            15'b00101110_0001_000: DATA = 1'b0;
            15'b00101110_0001_001: DATA = 1'b0;
            15'b00101110_0001_010: DATA = 1'b0;
            15'b00101110_0001_011: DATA = 1'b0;
            15'b00101110_0001_100: DATA = 1'b0;
            15'b00101110_0001_101: DATA = 1'b0;
            15'b00101110_0001_110: DATA = 1'b0;
            15'b00101110_0001_111: DATA = 1'b0;
            // . Row 2
            15'b00101110_0010_000: DATA = 1'b0;
            15'b00101110_0010_001: DATA = 1'b0;
            15'b00101110_0010_010: DATA = 1'b0;
            15'b00101110_0010_011: DATA = 1'b0;
            15'b00101110_0010_100: DATA = 1'b0;
            15'b00101110_0010_101: DATA = 1'b0;
            15'b00101110_0010_110: DATA = 1'b0;
            15'b00101110_0010_111: DATA = 1'b0;
            // . Row 3
            15'b00101110_0011_000: DATA = 1'b0;
            15'b00101110_0011_001: DATA = 1'b0;
            15'b00101110_0011_010: DATA = 1'b0;
            15'b00101110_0011_011: DATA = 1'b0;
            15'b00101110_0011_100: DATA = 1'b0;
            15'b00101110_0011_101: DATA = 1'b0;
            15'b00101110_0011_110: DATA = 1'b0;
            15'b00101110_0011_111: DATA = 1'b0;
            // . Row 4
            15'b00101110_0100_000: DATA = 1'b0;
            15'b00101110_0100_001: DATA = 1'b0;
            15'b00101110_0100_010: DATA = 1'b0;
            15'b00101110_0100_011: DATA = 1'b0;
            15'b00101110_0100_100: DATA = 1'b0;
            15'b00101110_0100_101: DATA = 1'b0;
            15'b00101110_0100_110: DATA = 1'b0;
            15'b00101110_0100_111: DATA = 1'b0;
            // . Row 5
            15'b00101110_0101_000: DATA = 1'b0;
            15'b00101110_0101_001: DATA = 1'b0;
            15'b00101110_0101_010: DATA = 1'b0;
            15'b00101110_0101_011: DATA = 1'b0;
            15'b00101110_0101_100: DATA = 1'b0;
            15'b00101110_0101_101: DATA = 1'b0;
            15'b00101110_0101_110: DATA = 1'b0;
            15'b00101110_0101_111: DATA = 1'b0;
            // . Row 6
            15'b00101110_0110_000: DATA = 1'b0;
            15'b00101110_0110_001: DATA = 1'b0;
            15'b00101110_0110_010: DATA = 1'b0;
            15'b00101110_0110_011: DATA = 1'b0;
            15'b00101110_0110_100: DATA = 1'b0;
            15'b00101110_0110_101: DATA = 1'b0;
            15'b00101110_0110_110: DATA = 1'b0;
            15'b00101110_0110_111: DATA = 1'b0;
            // . Row 7
            15'b00101110_0111_000: DATA = 1'b0;
            15'b00101110_0111_001: DATA = 1'b0;
            15'b00101110_0111_010: DATA = 1'b0;
            15'b00101110_0111_011: DATA = 1'b0;
            15'b00101110_0111_100: DATA = 1'b0;
            15'b00101110_0111_101: DATA = 1'b0;
            15'b00101110_0111_110: DATA = 1'b0;
            15'b00101110_0111_111: DATA = 1'b0;
            // . Row 8
            15'b00101110_1000_000: DATA = 1'b0;
            15'b00101110_1000_001: DATA = 1'b0;
            15'b00101110_1000_010: DATA = 1'b0;
            15'b00101110_1000_011: DATA = 1'b0;
            15'b00101110_1000_100: DATA = 1'b0;
            15'b00101110_1000_101: DATA = 1'b0;
            15'b00101110_1000_110: DATA = 1'b0;
            15'b00101110_1000_111: DATA = 1'b0;
            // . Row 9
            15'b00101110_1001_000: DATA = 1'b0;
            15'b00101110_1001_001: DATA = 1'b0;
            15'b00101110_1001_010: DATA = 1'b0;
            15'b00101110_1001_011: DATA = 1'b0;
            15'b00101110_1001_100: DATA = 1'b0;
            15'b00101110_1001_101: DATA = 1'b0;
            15'b00101110_1001_110: DATA = 1'b0;
            15'b00101110_1001_111: DATA = 1'b0;
            // . Row 10
            15'b00101110_1010_000: DATA = 1'b0;
            15'b00101110_1010_001: DATA = 1'b0;
            15'b00101110_1010_010: DATA = 1'b0;
            15'b00101110_1010_011: DATA = 1'b0;
            15'b00101110_1010_100: DATA = 1'b0;
            15'b00101110_1010_101: DATA = 1'b0;
            15'b00101110_1010_110: DATA = 1'b0;
            15'b00101110_1010_111: DATA = 1'b0;
            // . Row 11
            15'b00101110_1011_000: DATA = 1'b0;
            15'b00101110_1011_001: DATA = 1'b1;
            15'b00101110_1011_010: DATA = 1'b1;
            15'b00101110_1011_011: DATA = 1'b0;
            15'b00101110_1011_100: DATA = 1'b0;
            15'b00101110_1011_101: DATA = 1'b0;
            15'b00101110_1011_110: DATA = 1'b0;
            15'b00101110_1011_111: DATA = 1'b0;
            // . Row 12
            15'b00101110_1100_000: DATA = 1'b0;
            15'b00101110_1100_001: DATA = 1'b1;
            15'b00101110_1100_010: DATA = 1'b1;
            15'b00101110_1100_011: DATA = 1'b0;
            15'b00101110_1100_100: DATA = 1'b0;
            15'b00101110_1100_101: DATA = 1'b0;
            15'b00101110_1100_110: DATA = 1'b0;
            15'b00101110_1100_111: DATA = 1'b0;
            // . Row 13
            15'b00101110_1101_000: DATA = 1'b0;
            15'b00101110_1101_001: DATA = 1'b0;
            15'b00101110_1101_010: DATA = 1'b0;
            15'b00101110_1101_011: DATA = 1'b0;
            15'b00101110_1101_100: DATA = 1'b0;
            15'b00101110_1101_101: DATA = 1'b0;
            15'b00101110_1101_110: DATA = 1'b0;
            15'b00101110_1101_111: DATA = 1'b0;
            // . Row 14
            15'b00101110_1110_000: DATA = 1'b0;
            15'b00101110_1110_001: DATA = 1'b0;
            15'b00101110_1110_010: DATA = 1'b0;
            15'b00101110_1110_011: DATA = 1'b0;
            15'b00101110_1110_100: DATA = 1'b0;
            15'b00101110_1110_101: DATA = 1'b0;
            15'b00101110_1110_110: DATA = 1'b0;
            15'b00101110_1110_111: DATA = 1'b0;
            // . Row 15
            15'b00101110_1111_000: DATA = 1'b0;
            15'b00101110_1111_001: DATA = 1'b0;
            15'b00101110_1111_010: DATA = 1'b0;
            15'b00101110_1111_011: DATA = 1'b0;
            15'b00101110_1111_100: DATA = 1'b0;
            15'b00101110_1111_101: DATA = 1'b0;
            15'b00101110_1111_110: DATA = 1'b0;
            15'b00101110_1111_111: DATA = 1'b0;
            // 0 Row 0
            15'b00110000_0000_000: DATA = 1'b0;
            15'b00110000_0000_001: DATA = 1'b0;
            15'b00110000_0000_010: DATA = 1'b0;
            15'b00110000_0000_011: DATA = 1'b0;
            15'b00110000_0000_100: DATA = 1'b0;
            15'b00110000_0000_101: DATA = 1'b0;
            15'b00110000_0000_110: DATA = 1'b0;
            15'b00110000_0000_111: DATA = 1'b0;
            // 0 Row 1
            15'b00110000_0001_000: DATA = 1'b0;
            15'b00110000_0001_001: DATA = 1'b0;
            15'b00110000_0001_010: DATA = 1'b0;
            15'b00110000_0001_011: DATA = 1'b0;
            15'b00110000_0001_100: DATA = 1'b0;
            15'b00110000_0001_101: DATA = 1'b0;
            15'b00110000_0001_110: DATA = 1'b0;
            15'b00110000_0001_111: DATA = 1'b0;
            // 0 Row 2
            15'b00110000_0010_000: DATA = 1'b0;
            15'b00110000_0010_001: DATA = 1'b0;
            15'b00110000_0010_010: DATA = 1'b0;
            15'b00110000_0010_011: DATA = 1'b0;
            15'b00110000_0010_100: DATA = 1'b0;
            15'b00110000_0010_101: DATA = 1'b0;
            15'b00110000_0010_110: DATA = 1'b0;
            15'b00110000_0010_111: DATA = 1'b0;
            // 0 Row 3
            15'b00110000_0011_000: DATA = 1'b0;
            15'b00110000_0011_001: DATA = 1'b0;
            15'b00110000_0011_010: DATA = 1'b1;
            15'b00110000_0011_011: DATA = 1'b1;
            15'b00110000_0011_100: DATA = 1'b1;
            15'b00110000_0011_101: DATA = 1'b0;
            15'b00110000_0011_110: DATA = 1'b0;
            15'b00110000_0011_111: DATA = 1'b0;
            // 0 Row 4
            15'b00110000_0100_000: DATA = 1'b0;
            15'b00110000_0100_001: DATA = 1'b1;
            15'b00110000_0100_010: DATA = 1'b1;
            15'b00110000_0100_011: DATA = 1'b1;
            15'b00110000_0100_100: DATA = 1'b1;
            15'b00110000_0100_101: DATA = 1'b1;
            15'b00110000_0100_110: DATA = 1'b0;
            15'b00110000_0100_111: DATA = 1'b0;
            // 0 Row 5
            15'b00110000_0101_000: DATA = 1'b1;
            15'b00110000_0101_001: DATA = 1'b1;
            15'b00110000_0101_010: DATA = 1'b1;
            15'b00110000_0101_011: DATA = 1'b0;
            15'b00110000_0101_100: DATA = 1'b0;
            15'b00110000_0101_101: DATA = 1'b1;
            15'b00110000_0101_110: DATA = 1'b1;
            15'b00110000_0101_111: DATA = 1'b0;
            // 0 Row 6
            15'b00110000_0110_000: DATA = 1'b1;
            15'b00110000_0110_001: DATA = 1'b1;
            15'b00110000_0110_010: DATA = 1'b1;
            15'b00110000_0110_011: DATA = 1'b1;
            15'b00110000_0110_100: DATA = 1'b0;
            15'b00110000_0110_101: DATA = 1'b1;
            15'b00110000_0110_110: DATA = 1'b1;
            15'b00110000_0110_111: DATA = 1'b0;
            // 0 Row 7
            15'b00110000_0111_000: DATA = 1'b1;
            15'b00110000_0111_001: DATA = 1'b1;
            15'b00110000_0111_010: DATA = 1'b0;
            15'b00110000_0111_011: DATA = 1'b1;
            15'b00110000_0111_100: DATA = 1'b0;
            15'b00110000_0111_101: DATA = 1'b1;
            15'b00110000_0111_110: DATA = 1'b1;
            15'b00110000_0111_111: DATA = 1'b0;
            // 0 Row 8
            15'b00110000_1000_000: DATA = 1'b1;
            15'b00110000_1000_001: DATA = 1'b1;
            15'b00110000_1000_010: DATA = 1'b0;
            15'b00110000_1000_011: DATA = 1'b1;
            15'b00110000_1000_100: DATA = 1'b0;
            15'b00110000_1000_101: DATA = 1'b1;
            15'b00110000_1000_110: DATA = 1'b1;
            15'b00110000_1000_111: DATA = 1'b0;
            // 0 Row 9
            15'b00110000_1001_000: DATA = 1'b1;
            15'b00110000_1001_001: DATA = 1'b1;
            15'b00110000_1001_010: DATA = 1'b0;
            15'b00110000_1001_011: DATA = 1'b1;
            15'b00110000_1001_100: DATA = 1'b1;
            15'b00110000_1001_101: DATA = 1'b1;
            15'b00110000_1001_110: DATA = 1'b1;
            15'b00110000_1001_111: DATA = 1'b0;
            // 0 Row 10
            15'b00110000_1010_000: DATA = 1'b1;
            15'b00110000_1010_001: DATA = 1'b1;
            15'b00110000_1010_010: DATA = 1'b0;
            15'b00110000_1010_011: DATA = 1'b0;
            15'b00110000_1010_100: DATA = 1'b1;
            15'b00110000_1010_101: DATA = 1'b1;
            15'b00110000_1010_110: DATA = 1'b1;
            15'b00110000_1010_111: DATA = 1'b0;
            // 0 Row 11
            15'b00110000_1011_000: DATA = 1'b0;
            15'b00110000_1011_001: DATA = 1'b1;
            15'b00110000_1011_010: DATA = 1'b1;
            15'b00110000_1011_011: DATA = 1'b1;
            15'b00110000_1011_100: DATA = 1'b1;
            15'b00110000_1011_101: DATA = 1'b1;
            15'b00110000_1011_110: DATA = 1'b0;
            15'b00110000_1011_111: DATA = 1'b0;
            // 0 Row 12
            15'b00110000_1100_000: DATA = 1'b0;
            15'b00110000_1100_001: DATA = 1'b0;
            15'b00110000_1100_010: DATA = 1'b1;
            15'b00110000_1100_011: DATA = 1'b1;
            15'b00110000_1100_100: DATA = 1'b1;
            15'b00110000_1100_101: DATA = 1'b0;
            15'b00110000_1100_110: DATA = 1'b0;
            15'b00110000_1100_111: DATA = 1'b0;
            // 0 Row 13
            15'b00110000_1101_000: DATA = 1'b0;
            15'b00110000_1101_001: DATA = 1'b0;
            15'b00110000_1101_010: DATA = 1'b0;
            15'b00110000_1101_011: DATA = 1'b0;
            15'b00110000_1101_100: DATA = 1'b0;
            15'b00110000_1101_101: DATA = 1'b0;
            15'b00110000_1101_110: DATA = 1'b0;
            15'b00110000_1101_111: DATA = 1'b0;
            // 0 Row 14
            15'b00110000_1110_000: DATA = 1'b0;
            15'b00110000_1110_001: DATA = 1'b0;
            15'b00110000_1110_010: DATA = 1'b0;
            15'b00110000_1110_011: DATA = 1'b0;
            15'b00110000_1110_100: DATA = 1'b0;
            15'b00110000_1110_101: DATA = 1'b0;
            15'b00110000_1110_110: DATA = 1'b0;
            15'b00110000_1110_111: DATA = 1'b0;
            // 0 Row 15
            15'b00110000_1111_000: DATA = 1'b0;
            15'b00110000_1111_001: DATA = 1'b0;
            15'b00110000_1111_010: DATA = 1'b0;
            15'b00110000_1111_011: DATA = 1'b0;
            15'b00110000_1111_100: DATA = 1'b0;
            15'b00110000_1111_101: DATA = 1'b0;
            15'b00110000_1111_110: DATA = 1'b0;
            15'b00110000_1111_111: DATA = 1'b0;
            // 1 Row 0
            15'b00110001_0000_000: DATA = 1'b0;
            15'b00110001_0000_001: DATA = 1'b0;
            15'b00110001_0000_010: DATA = 1'b0;
            15'b00110001_0000_011: DATA = 1'b0;
            15'b00110001_0000_100: DATA = 1'b0;
            15'b00110001_0000_101: DATA = 1'b0;
            15'b00110001_0000_110: DATA = 1'b0;
            15'b00110001_0000_111: DATA = 1'b0;
            // 1 Row 1
            15'b00110001_0001_000: DATA = 1'b0;
            15'b00110001_0001_001: DATA = 1'b0;
            15'b00110001_0001_010: DATA = 1'b0;
            15'b00110001_0001_011: DATA = 1'b0;
            15'b00110001_0001_100: DATA = 1'b0;
            15'b00110001_0001_101: DATA = 1'b0;
            15'b00110001_0001_110: DATA = 1'b0;
            15'b00110001_0001_111: DATA = 1'b0;
            // 1 Row 2
            15'b00110001_0010_000: DATA = 1'b0;
            15'b00110001_0010_001: DATA = 1'b0;
            15'b00110001_0010_010: DATA = 1'b0;
            15'b00110001_0010_011: DATA = 1'b0;
            15'b00110001_0010_100: DATA = 1'b0;
            15'b00110001_0010_101: DATA = 1'b0;
            15'b00110001_0010_110: DATA = 1'b0;
            15'b00110001_0010_111: DATA = 1'b0;
            // 1 Row 3
            15'b00110001_0011_000: DATA = 1'b0;
            15'b00110001_0011_001: DATA = 1'b0;
            15'b00110001_0011_010: DATA = 1'b1;
            15'b00110001_0011_011: DATA = 1'b1;
            15'b00110001_0011_100: DATA = 1'b1;
            15'b00110001_0011_101: DATA = 1'b0;
            15'b00110001_0011_110: DATA = 1'b0;
            15'b00110001_0011_111: DATA = 1'b0;
            // 1 Row 4
            15'b00110001_0100_000: DATA = 1'b0;
            15'b00110001_0100_001: DATA = 1'b1;
            15'b00110001_0100_010: DATA = 1'b1;
            15'b00110001_0100_011: DATA = 1'b1;
            15'b00110001_0100_100: DATA = 1'b1;
            15'b00110001_0100_101: DATA = 1'b0;
            15'b00110001_0100_110: DATA = 1'b0;
            15'b00110001_0100_111: DATA = 1'b0;
            // 1 Row 5
            15'b00110001_0101_000: DATA = 1'b1;
            15'b00110001_0101_001: DATA = 1'b1;
            15'b00110001_0101_010: DATA = 1'b0;
            15'b00110001_0101_011: DATA = 1'b1;
            15'b00110001_0101_100: DATA = 1'b1;
            15'b00110001_0101_101: DATA = 1'b0;
            15'b00110001_0101_110: DATA = 1'b0;
            15'b00110001_0101_111: DATA = 1'b0;
            // 1 Row 6
            15'b00110001_0110_000: DATA = 1'b0;
            15'b00110001_0110_001: DATA = 1'b0;
            15'b00110001_0110_010: DATA = 1'b0;
            15'b00110001_0110_011: DATA = 1'b1;
            15'b00110001_0110_100: DATA = 1'b1;
            15'b00110001_0110_101: DATA = 1'b0;
            15'b00110001_0110_110: DATA = 1'b0;
            15'b00110001_0110_111: DATA = 1'b0;
            // 1 Row 7
            15'b00110001_0111_000: DATA = 1'b0;
            15'b00110001_0111_001: DATA = 1'b0;
            15'b00110001_0111_010: DATA = 1'b0;
            15'b00110001_0111_011: DATA = 1'b1;
            15'b00110001_0111_100: DATA = 1'b1;
            15'b00110001_0111_101: DATA = 1'b0;
            15'b00110001_0111_110: DATA = 1'b0;
            15'b00110001_0111_111: DATA = 1'b0;
            // 1 Row 8
            15'b00110001_1000_000: DATA = 1'b0;
            15'b00110001_1000_001: DATA = 1'b0;
            15'b00110001_1000_010: DATA = 1'b0;
            15'b00110001_1000_011: DATA = 1'b1;
            15'b00110001_1000_100: DATA = 1'b1;
            15'b00110001_1000_101: DATA = 1'b0;
            15'b00110001_1000_110: DATA = 1'b0;
            15'b00110001_1000_111: DATA = 1'b0;
            // 1 Row 9
            15'b00110001_1001_000: DATA = 1'b0;
            15'b00110001_1001_001: DATA = 1'b0;
            15'b00110001_1001_010: DATA = 1'b0;
            15'b00110001_1001_011: DATA = 1'b1;
            15'b00110001_1001_100: DATA = 1'b1;
            15'b00110001_1001_101: DATA = 1'b0;
            15'b00110001_1001_110: DATA = 1'b0;
            15'b00110001_1001_111: DATA = 1'b0;
            // 1 Row 10
            15'b00110001_1010_000: DATA = 1'b0;
            15'b00110001_1010_001: DATA = 1'b0;
            15'b00110001_1010_010: DATA = 1'b0;
            15'b00110001_1010_011: DATA = 1'b1;
            15'b00110001_1010_100: DATA = 1'b1;
            15'b00110001_1010_101: DATA = 1'b0;
            15'b00110001_1010_110: DATA = 1'b0;
            15'b00110001_1010_111: DATA = 1'b0;
            // 1 Row 11
            15'b00110001_1011_000: DATA = 1'b1;
            15'b00110001_1011_001: DATA = 1'b1;
            15'b00110001_1011_010: DATA = 1'b1;
            15'b00110001_1011_011: DATA = 1'b1;
            15'b00110001_1011_100: DATA = 1'b1;
            15'b00110001_1011_101: DATA = 1'b1;
            15'b00110001_1011_110: DATA = 1'b1;
            15'b00110001_1011_111: DATA = 1'b0;
            // 1 Row 12
            15'b00110001_1100_000: DATA = 1'b1;
            15'b00110001_1100_001: DATA = 1'b1;
            15'b00110001_1100_010: DATA = 1'b1;
            15'b00110001_1100_011: DATA = 1'b1;
            15'b00110001_1100_100: DATA = 1'b1;
            15'b00110001_1100_101: DATA = 1'b1;
            15'b00110001_1100_110: DATA = 1'b1;
            15'b00110001_1100_111: DATA = 1'b0;
            // 1 Row 13
            15'b00110001_1101_000: DATA = 1'b0;
            15'b00110001_1101_001: DATA = 1'b0;
            15'b00110001_1101_010: DATA = 1'b0;
            15'b00110001_1101_011: DATA = 1'b0;
            15'b00110001_1101_100: DATA = 1'b0;
            15'b00110001_1101_101: DATA = 1'b0;
            15'b00110001_1101_110: DATA = 1'b0;
            15'b00110001_1101_111: DATA = 1'b0;
            // 1 Row 14
            15'b00110001_1110_000: DATA = 1'b0;
            15'b00110001_1110_001: DATA = 1'b0;
            15'b00110001_1110_010: DATA = 1'b0;
            15'b00110001_1110_011: DATA = 1'b0;
            15'b00110001_1110_100: DATA = 1'b0;
            15'b00110001_1110_101: DATA = 1'b0;
            15'b00110001_1110_110: DATA = 1'b0;
            15'b00110001_1110_111: DATA = 1'b0;
            // 1 Row 15
            15'b00110001_1111_000: DATA = 1'b0;
            15'b00110001_1111_001: DATA = 1'b0;
            15'b00110001_1111_010: DATA = 1'b0;
            15'b00110001_1111_011: DATA = 1'b0;
            15'b00110001_1111_100: DATA = 1'b0;
            15'b00110001_1111_101: DATA = 1'b0;
            15'b00110001_1111_110: DATA = 1'b0;
            15'b00110001_1111_111: DATA = 1'b0;
            // 2 Row 0
            15'b00110010_0000_000: DATA = 1'b0;
            15'b00110010_0000_001: DATA = 1'b0;
            15'b00110010_0000_010: DATA = 1'b0;
            15'b00110010_0000_011: DATA = 1'b0;
            15'b00110010_0000_100: DATA = 1'b0;
            15'b00110010_0000_101: DATA = 1'b0;
            15'b00110010_0000_110: DATA = 1'b0;
            15'b00110010_0000_111: DATA = 1'b0;
            // 2 Row 1
            15'b00110010_0001_000: DATA = 1'b0;
            15'b00110010_0001_001: DATA = 1'b0;
            15'b00110010_0001_010: DATA = 1'b0;
            15'b00110010_0001_011: DATA = 1'b0;
            15'b00110010_0001_100: DATA = 1'b0;
            15'b00110010_0001_101: DATA = 1'b0;
            15'b00110010_0001_110: DATA = 1'b0;
            15'b00110010_0001_111: DATA = 1'b0;
            // 2 Row 2
            15'b00110010_0010_000: DATA = 1'b0;
            15'b00110010_0010_001: DATA = 1'b0;
            15'b00110010_0010_010: DATA = 1'b0;
            15'b00110010_0010_011: DATA = 1'b0;
            15'b00110010_0010_100: DATA = 1'b0;
            15'b00110010_0010_101: DATA = 1'b0;
            15'b00110010_0010_110: DATA = 1'b0;
            15'b00110010_0010_111: DATA = 1'b0;
            // 2 Row 3
            15'b00110010_0011_000: DATA = 1'b0;
            15'b00110010_0011_001: DATA = 1'b0;
            15'b00110010_0011_010: DATA = 1'b1;
            15'b00110010_0011_011: DATA = 1'b1;
            15'b00110010_0011_100: DATA = 1'b1;
            15'b00110010_0011_101: DATA = 1'b0;
            15'b00110010_0011_110: DATA = 1'b0;
            15'b00110010_0011_111: DATA = 1'b0;
            // 2 Row 4
            15'b00110010_0100_000: DATA = 1'b0;
            15'b00110010_0100_001: DATA = 1'b1;
            15'b00110010_0100_010: DATA = 1'b1;
            15'b00110010_0100_011: DATA = 1'b0;
            15'b00110010_0100_100: DATA = 1'b1;
            15'b00110010_0100_101: DATA = 1'b1;
            15'b00110010_0100_110: DATA = 1'b0;
            15'b00110010_0100_111: DATA = 1'b0;
            // 2 Row 5
            15'b00110010_0101_000: DATA = 1'b1;
            15'b00110010_0101_001: DATA = 1'b1;
            15'b00110010_0101_010: DATA = 1'b0;
            15'b00110010_0101_011: DATA = 1'b0;
            15'b00110010_0101_100: DATA = 1'b0;
            15'b00110010_0101_101: DATA = 1'b1;
            15'b00110010_0101_110: DATA = 1'b1;
            15'b00110010_0101_111: DATA = 1'b0;
            // 2 Row 6
            15'b00110010_0110_000: DATA = 1'b0;
            15'b00110010_0110_001: DATA = 1'b0;
            15'b00110010_0110_010: DATA = 1'b0;
            15'b00110010_0110_011: DATA = 1'b0;
            15'b00110010_0110_100: DATA = 1'b0;
            15'b00110010_0110_101: DATA = 1'b1;
            15'b00110010_0110_110: DATA = 1'b1;
            15'b00110010_0110_111: DATA = 1'b0;
            // 2 Row 7
            15'b00110010_0111_000: DATA = 1'b0;
            15'b00110010_0111_001: DATA = 1'b0;
            15'b00110010_0111_010: DATA = 1'b0;
            15'b00110010_0111_011: DATA = 1'b0;
            15'b00110010_0111_100: DATA = 1'b1;
            15'b00110010_0111_101: DATA = 1'b1;
            15'b00110010_0111_110: DATA = 1'b0;
            15'b00110010_0111_111: DATA = 1'b0;
            // 2 Row 8
            15'b00110010_1000_000: DATA = 1'b0;
            15'b00110010_1000_001: DATA = 1'b0;
            15'b00110010_1000_010: DATA = 1'b0;
            15'b00110010_1000_011: DATA = 1'b1;
            15'b00110010_1000_100: DATA = 1'b1;
            15'b00110010_1000_101: DATA = 1'b0;
            15'b00110010_1000_110: DATA = 1'b0;
            15'b00110010_1000_111: DATA = 1'b0;
            // 2 Row 9
            15'b00110010_1001_000: DATA = 1'b0;
            15'b00110010_1001_001: DATA = 1'b0;
            15'b00110010_1001_010: DATA = 1'b1;
            15'b00110010_1001_011: DATA = 1'b1;
            15'b00110010_1001_100: DATA = 1'b0;
            15'b00110010_1001_101: DATA = 1'b0;
            15'b00110010_1001_110: DATA = 1'b0;
            15'b00110010_1001_111: DATA = 1'b0;
            // 2 Row 10
            15'b00110010_1010_000: DATA = 1'b0;
            15'b00110010_1010_001: DATA = 1'b1;
            15'b00110010_1010_010: DATA = 1'b1;
            15'b00110010_1010_011: DATA = 1'b0;
            15'b00110010_1010_100: DATA = 1'b0;
            15'b00110010_1010_101: DATA = 1'b0;
            15'b00110010_1010_110: DATA = 1'b0;
            15'b00110010_1010_111: DATA = 1'b0;
            // 2 Row 11
            15'b00110010_1011_000: DATA = 1'b1;
            15'b00110010_1011_001: DATA = 1'b1;
            15'b00110010_1011_010: DATA = 1'b1;
            15'b00110010_1011_011: DATA = 1'b1;
            15'b00110010_1011_100: DATA = 1'b1;
            15'b00110010_1011_101: DATA = 1'b1;
            15'b00110010_1011_110: DATA = 1'b1;
            15'b00110010_1011_111: DATA = 1'b0;
            // 2 Row 12
            15'b00110010_1100_000: DATA = 1'b1;
            15'b00110010_1100_001: DATA = 1'b1;
            15'b00110010_1100_010: DATA = 1'b1;
            15'b00110010_1100_011: DATA = 1'b1;
            15'b00110010_1100_100: DATA = 1'b1;
            15'b00110010_1100_101: DATA = 1'b1;
            15'b00110010_1100_110: DATA = 1'b1;
            15'b00110010_1100_111: DATA = 1'b0;
            // 2 Row 13
            15'b00110010_1101_000: DATA = 1'b0;
            15'b00110010_1101_001: DATA = 1'b0;
            15'b00110010_1101_010: DATA = 1'b0;
            15'b00110010_1101_011: DATA = 1'b0;
            15'b00110010_1101_100: DATA = 1'b0;
            15'b00110010_1101_101: DATA = 1'b0;
            15'b00110010_1101_110: DATA = 1'b0;
            15'b00110010_1101_111: DATA = 1'b0;
            // 2 Row 14
            15'b00110010_1110_000: DATA = 1'b0;
            15'b00110010_1110_001: DATA = 1'b0;
            15'b00110010_1110_010: DATA = 1'b0;
            15'b00110010_1110_011: DATA = 1'b0;
            15'b00110010_1110_100: DATA = 1'b0;
            15'b00110010_1110_101: DATA = 1'b0;
            15'b00110010_1110_110: DATA = 1'b0;
            15'b00110010_1110_111: DATA = 1'b0;
            // 2 Row 15
            15'b00110010_1111_000: DATA = 1'b0;
            15'b00110010_1111_001: DATA = 1'b0;
            15'b00110010_1111_010: DATA = 1'b0;
            15'b00110010_1111_011: DATA = 1'b0;
            15'b00110010_1111_100: DATA = 1'b0;
            15'b00110010_1111_101: DATA = 1'b0;
            15'b00110010_1111_110: DATA = 1'b0;
            15'b00110010_1111_111: DATA = 1'b0;
            // 3 Row 0
            15'b00110011_0000_000: DATA = 1'b0;
            15'b00110011_0000_001: DATA = 1'b0;
            15'b00110011_0000_010: DATA = 1'b0;
            15'b00110011_0000_011: DATA = 1'b0;
            15'b00110011_0000_100: DATA = 1'b0;
            15'b00110011_0000_101: DATA = 1'b0;
            15'b00110011_0000_110: DATA = 1'b0;
            15'b00110011_0000_111: DATA = 1'b0;
            // 3 Row 1
            15'b00110011_0001_000: DATA = 1'b0;
            15'b00110011_0001_001: DATA = 1'b0;
            15'b00110011_0001_010: DATA = 1'b0;
            15'b00110011_0001_011: DATA = 1'b0;
            15'b00110011_0001_100: DATA = 1'b0;
            15'b00110011_0001_101: DATA = 1'b0;
            15'b00110011_0001_110: DATA = 1'b0;
            15'b00110011_0001_111: DATA = 1'b0;
            // 3 Row 2
            15'b00110011_0010_000: DATA = 1'b0;
            15'b00110011_0010_001: DATA = 1'b0;
            15'b00110011_0010_010: DATA = 1'b0;
            15'b00110011_0010_011: DATA = 1'b0;
            15'b00110011_0010_100: DATA = 1'b0;
            15'b00110011_0010_101: DATA = 1'b0;
            15'b00110011_0010_110: DATA = 1'b0;
            15'b00110011_0010_111: DATA = 1'b0;
            // 3 Row 3
            15'b00110011_0011_000: DATA = 1'b0;
            15'b00110011_0011_001: DATA = 1'b0;
            15'b00110011_0011_010: DATA = 1'b1;
            15'b00110011_0011_011: DATA = 1'b1;
            15'b00110011_0011_100: DATA = 1'b1;
            15'b00110011_0011_101: DATA = 1'b0;
            15'b00110011_0011_110: DATA = 1'b0;
            15'b00110011_0011_111: DATA = 1'b0;
            // 3 Row 4
            15'b00110011_0100_000: DATA = 1'b0;
            15'b00110011_0100_001: DATA = 1'b1;
            15'b00110011_0100_010: DATA = 1'b1;
            15'b00110011_0100_011: DATA = 1'b0;
            15'b00110011_0100_100: DATA = 1'b1;
            15'b00110011_0100_101: DATA = 1'b1;
            15'b00110011_0100_110: DATA = 1'b0;
            15'b00110011_0100_111: DATA = 1'b0;
            // 3 Row 5
            15'b00110011_0101_000: DATA = 1'b1;
            15'b00110011_0101_001: DATA = 1'b1;
            15'b00110011_0101_010: DATA = 1'b0;
            15'b00110011_0101_011: DATA = 1'b0;
            15'b00110011_0101_100: DATA = 1'b0;
            15'b00110011_0101_101: DATA = 1'b1;
            15'b00110011_0101_110: DATA = 1'b1;
            15'b00110011_0101_111: DATA = 1'b0;
            // 3 Row 6
            15'b00110011_0110_000: DATA = 1'b0;
            15'b00110011_0110_001: DATA = 1'b0;
            15'b00110011_0110_010: DATA = 1'b0;
            15'b00110011_0110_011: DATA = 1'b0;
            15'b00110011_0110_100: DATA = 1'b0;
            15'b00110011_0110_101: DATA = 1'b1;
            15'b00110011_0110_110: DATA = 1'b1;
            15'b00110011_0110_111: DATA = 1'b0;
            // 3 Row 7
            15'b00110011_0111_000: DATA = 1'b0;
            15'b00110011_0111_001: DATA = 1'b0;
            15'b00110011_0111_010: DATA = 1'b0;
            15'b00110011_0111_011: DATA = 1'b1;
            15'b00110011_0111_100: DATA = 1'b1;
            15'b00110011_0111_101: DATA = 1'b1;
            15'b00110011_0111_110: DATA = 1'b0;
            15'b00110011_0111_111: DATA = 1'b0;
            // 3 Row 8
            15'b00110011_1000_000: DATA = 1'b0;
            15'b00110011_1000_001: DATA = 1'b0;
            15'b00110011_1000_010: DATA = 1'b0;
            15'b00110011_1000_011: DATA = 1'b1;
            15'b00110011_1000_100: DATA = 1'b1;
            15'b00110011_1000_101: DATA = 1'b1;
            15'b00110011_1000_110: DATA = 1'b0;
            15'b00110011_1000_111: DATA = 1'b0;
            // 3 Row 9
            15'b00110011_1001_000: DATA = 1'b0;
            15'b00110011_1001_001: DATA = 1'b0;
            15'b00110011_1001_010: DATA = 1'b0;
            15'b00110011_1001_011: DATA = 1'b0;
            15'b00110011_1001_100: DATA = 1'b0;
            15'b00110011_1001_101: DATA = 1'b1;
            15'b00110011_1001_110: DATA = 1'b1;
            15'b00110011_1001_111: DATA = 1'b0;
            // 3 Row 10
            15'b00110011_1010_000: DATA = 1'b1;
            15'b00110011_1010_001: DATA = 1'b1;
            15'b00110011_1010_010: DATA = 1'b0;
            15'b00110011_1010_011: DATA = 1'b0;
            15'b00110011_1010_100: DATA = 1'b0;
            15'b00110011_1010_101: DATA = 1'b1;
            15'b00110011_1010_110: DATA = 1'b1;
            15'b00110011_1010_111: DATA = 1'b0;
            // 3 Row 11
            15'b00110011_1011_000: DATA = 1'b0;
            15'b00110011_1011_001: DATA = 1'b1;
            15'b00110011_1011_010: DATA = 1'b1;
            15'b00110011_1011_011: DATA = 1'b0;
            15'b00110011_1011_100: DATA = 1'b1;
            15'b00110011_1011_101: DATA = 1'b1;
            15'b00110011_1011_110: DATA = 1'b0;
            15'b00110011_1011_111: DATA = 1'b0;
            // 3 Row 12
            15'b00110011_1100_000: DATA = 1'b0;
            15'b00110011_1100_001: DATA = 1'b0;
            15'b00110011_1100_010: DATA = 1'b1;
            15'b00110011_1100_011: DATA = 1'b1;
            15'b00110011_1100_100: DATA = 1'b1;
            15'b00110011_1100_101: DATA = 1'b0;
            15'b00110011_1100_110: DATA = 1'b0;
            15'b00110011_1100_111: DATA = 1'b0;
            // 3 Row 13
            15'b00110011_1101_000: DATA = 1'b0;
            15'b00110011_1101_001: DATA = 1'b0;
            15'b00110011_1101_010: DATA = 1'b0;
            15'b00110011_1101_011: DATA = 1'b0;
            15'b00110011_1101_100: DATA = 1'b0;
            15'b00110011_1101_101: DATA = 1'b0;
            15'b00110011_1101_110: DATA = 1'b0;
            15'b00110011_1101_111: DATA = 1'b0;
            // 3 Row 14
            15'b00110011_1110_000: DATA = 1'b0;
            15'b00110011_1110_001: DATA = 1'b0;
            15'b00110011_1110_010: DATA = 1'b0;
            15'b00110011_1110_011: DATA = 1'b0;
            15'b00110011_1110_100: DATA = 1'b0;
            15'b00110011_1110_101: DATA = 1'b0;
            15'b00110011_1110_110: DATA = 1'b0;
            15'b00110011_1110_111: DATA = 1'b0;
            // 3 Row 15
            15'b00110011_1111_000: DATA = 1'b0;
            15'b00110011_1111_001: DATA = 1'b0;
            15'b00110011_1111_010: DATA = 1'b0;
            15'b00110011_1111_011: DATA = 1'b0;
            15'b00110011_1111_100: DATA = 1'b0;
            15'b00110011_1111_101: DATA = 1'b0;
            15'b00110011_1111_110: DATA = 1'b0;
            15'b00110011_1111_111: DATA = 1'b0;
            // 4 Row 0
            15'b00110100_0000_000: DATA = 1'b0;
            15'b00110100_0000_001: DATA = 1'b0;
            15'b00110100_0000_010: DATA = 1'b0;
            15'b00110100_0000_011: DATA = 1'b0;
            15'b00110100_0000_100: DATA = 1'b0;
            15'b00110100_0000_101: DATA = 1'b0;
            15'b00110100_0000_110: DATA = 1'b0;
            15'b00110100_0000_111: DATA = 1'b0;
            // 4 Row 1
            15'b00110100_0001_000: DATA = 1'b0;
            15'b00110100_0001_001: DATA = 1'b0;
            15'b00110100_0001_010: DATA = 1'b0;
            15'b00110100_0001_011: DATA = 1'b0;
            15'b00110100_0001_100: DATA = 1'b0;
            15'b00110100_0001_101: DATA = 1'b0;
            15'b00110100_0001_110: DATA = 1'b0;
            15'b00110100_0001_111: DATA = 1'b0;
            // 4 Row 2
            15'b00110100_0010_000: DATA = 1'b0;
            15'b00110100_0010_001: DATA = 1'b0;
            15'b00110100_0010_010: DATA = 1'b0;
            15'b00110100_0010_011: DATA = 1'b0;
            15'b00110100_0010_100: DATA = 1'b0;
            15'b00110100_0010_101: DATA = 1'b0;
            15'b00110100_0010_110: DATA = 1'b0;
            15'b00110100_0010_111: DATA = 1'b0;
            // 4 Row 3
            15'b00110100_0011_000: DATA = 1'b0;
            15'b00110100_0011_001: DATA = 1'b0;
            15'b00110100_0011_010: DATA = 1'b0;
            15'b00110100_0011_011: DATA = 1'b0;
            15'b00110100_0011_100: DATA = 1'b1;
            15'b00110100_0011_101: DATA = 1'b1;
            15'b00110100_0011_110: DATA = 1'b0;
            15'b00110100_0011_111: DATA = 1'b0;
            // 4 Row 4
            15'b00110100_0100_000: DATA = 1'b0;
            15'b00110100_0100_001: DATA = 1'b0;
            15'b00110100_0100_010: DATA = 1'b0;
            15'b00110100_0100_011: DATA = 1'b1;
            15'b00110100_0100_100: DATA = 1'b1;
            15'b00110100_0100_101: DATA = 1'b1;
            15'b00110100_0100_110: DATA = 1'b0;
            15'b00110100_0100_111: DATA = 1'b0;
            // 4 Row 5
            15'b00110100_0101_000: DATA = 1'b0;
            15'b00110100_0101_001: DATA = 1'b0;
            15'b00110100_0101_010: DATA = 1'b1;
            15'b00110100_0101_011: DATA = 1'b1;
            15'b00110100_0101_100: DATA = 1'b1;
            15'b00110100_0101_101: DATA = 1'b1;
            15'b00110100_0101_110: DATA = 1'b0;
            15'b00110100_0101_111: DATA = 1'b0;
            // 4 Row 6
            15'b00110100_0110_000: DATA = 1'b0;
            15'b00110100_0110_001: DATA = 1'b1;
            15'b00110100_0110_010: DATA = 1'b1;
            15'b00110100_0110_011: DATA = 1'b0;
            15'b00110100_0110_100: DATA = 1'b1;
            15'b00110100_0110_101: DATA = 1'b1;
            15'b00110100_0110_110: DATA = 1'b0;
            15'b00110100_0110_111: DATA = 1'b0;
            // 4 Row 7
            15'b00110100_0111_000: DATA = 1'b1;
            15'b00110100_0111_001: DATA = 1'b1;
            15'b00110100_0111_010: DATA = 1'b0;
            15'b00110100_0111_011: DATA = 1'b0;
            15'b00110100_0111_100: DATA = 1'b1;
            15'b00110100_0111_101: DATA = 1'b1;
            15'b00110100_0111_110: DATA = 1'b0;
            15'b00110100_0111_111: DATA = 1'b0;
            // 4 Row 8
            15'b00110100_1000_000: DATA = 1'b1;
            15'b00110100_1000_001: DATA = 1'b0;
            15'b00110100_1000_010: DATA = 1'b0;
            15'b00110100_1000_011: DATA = 1'b0;
            15'b00110100_1000_100: DATA = 1'b1;
            15'b00110100_1000_101: DATA = 1'b1;
            15'b00110100_1000_110: DATA = 1'b0;
            15'b00110100_1000_111: DATA = 1'b0;
            // 4 Row 9
            15'b00110100_1001_000: DATA = 1'b1;
            15'b00110100_1001_001: DATA = 1'b1;
            15'b00110100_1001_010: DATA = 1'b1;
            15'b00110100_1001_011: DATA = 1'b1;
            15'b00110100_1001_100: DATA = 1'b1;
            15'b00110100_1001_101: DATA = 1'b1;
            15'b00110100_1001_110: DATA = 1'b1;
            15'b00110100_1001_111: DATA = 1'b0;
            // 4 Row 10
            15'b00110100_1010_000: DATA = 1'b1;
            15'b00110100_1010_001: DATA = 1'b1;
            15'b00110100_1010_010: DATA = 1'b1;
            15'b00110100_1010_011: DATA = 1'b1;
            15'b00110100_1010_100: DATA = 1'b1;
            15'b00110100_1010_101: DATA = 1'b1;
            15'b00110100_1010_110: DATA = 1'b1;
            15'b00110100_1010_111: DATA = 1'b0;
            // 4 Row 11
            15'b00110100_1011_000: DATA = 1'b0;
            15'b00110100_1011_001: DATA = 1'b0;
            15'b00110100_1011_010: DATA = 1'b0;
            15'b00110100_1011_011: DATA = 1'b0;
            15'b00110100_1011_100: DATA = 1'b1;
            15'b00110100_1011_101: DATA = 1'b1;
            15'b00110100_1011_110: DATA = 1'b0;
            15'b00110100_1011_111: DATA = 1'b0;
            // 4 Row 12
            15'b00110100_1100_000: DATA = 1'b0;
            15'b00110100_1100_001: DATA = 1'b0;
            15'b00110100_1100_010: DATA = 1'b0;
            15'b00110100_1100_011: DATA = 1'b0;
            15'b00110100_1100_100: DATA = 1'b1;
            15'b00110100_1100_101: DATA = 1'b1;
            15'b00110100_1100_110: DATA = 1'b0;
            15'b00110100_1100_111: DATA = 1'b0;
            // 4 Row 13
            15'b00110100_1101_000: DATA = 1'b0;
            15'b00110100_1101_001: DATA = 1'b0;
            15'b00110100_1101_010: DATA = 1'b0;
            15'b00110100_1101_011: DATA = 1'b0;
            15'b00110100_1101_100: DATA = 1'b0;
            15'b00110100_1101_101: DATA = 1'b0;
            15'b00110100_1101_110: DATA = 1'b0;
            15'b00110100_1101_111: DATA = 1'b0;
            // 4 Row 14
            15'b00110100_1110_000: DATA = 1'b0;
            15'b00110100_1110_001: DATA = 1'b0;
            15'b00110100_1110_010: DATA = 1'b0;
            15'b00110100_1110_011: DATA = 1'b0;
            15'b00110100_1110_100: DATA = 1'b0;
            15'b00110100_1110_101: DATA = 1'b0;
            15'b00110100_1110_110: DATA = 1'b0;
            15'b00110100_1110_111: DATA = 1'b0;
            // 4 Row 15
            15'b00110100_1111_000: DATA = 1'b0;
            15'b00110100_1111_001: DATA = 1'b0;
            15'b00110100_1111_010: DATA = 1'b0;
            15'b00110100_1111_011: DATA = 1'b0;
            15'b00110100_1111_100: DATA = 1'b0;
            15'b00110100_1111_101: DATA = 1'b0;
            15'b00110100_1111_110: DATA = 1'b0;
            15'b00110100_1111_111: DATA = 1'b0;
            // 5 Row 0
            15'b00110101_0000_000: DATA = 1'b0;
            15'b00110101_0000_001: DATA = 1'b0;
            15'b00110101_0000_010: DATA = 1'b0;
            15'b00110101_0000_011: DATA = 1'b0;
            15'b00110101_0000_100: DATA = 1'b0;
            15'b00110101_0000_101: DATA = 1'b0;
            15'b00110101_0000_110: DATA = 1'b0;
            15'b00110101_0000_111: DATA = 1'b0;
            // 5 Row 1
            15'b00110101_0001_000: DATA = 1'b0;
            15'b00110101_0001_001: DATA = 1'b0;
            15'b00110101_0001_010: DATA = 1'b0;
            15'b00110101_0001_011: DATA = 1'b0;
            15'b00110101_0001_100: DATA = 1'b0;
            15'b00110101_0001_101: DATA = 1'b0;
            15'b00110101_0001_110: DATA = 1'b0;
            15'b00110101_0001_111: DATA = 1'b0;
            // 5 Row 2
            15'b00110101_0010_000: DATA = 1'b0;
            15'b00110101_0010_001: DATA = 1'b0;
            15'b00110101_0010_010: DATA = 1'b0;
            15'b00110101_0010_011: DATA = 1'b0;
            15'b00110101_0010_100: DATA = 1'b0;
            15'b00110101_0010_101: DATA = 1'b0;
            15'b00110101_0010_110: DATA = 1'b0;
            15'b00110101_0010_111: DATA = 1'b0;
            // 5 Row 3
            15'b00110101_0011_000: DATA = 1'b1;
            15'b00110101_0011_001: DATA = 1'b1;
            15'b00110101_0011_010: DATA = 1'b1;
            15'b00110101_0011_011: DATA = 1'b1;
            15'b00110101_0011_100: DATA = 1'b1;
            15'b00110101_0011_101: DATA = 1'b1;
            15'b00110101_0011_110: DATA = 1'b1;
            15'b00110101_0011_111: DATA = 1'b0;
            // 5 Row 4
            15'b00110101_0100_000: DATA = 1'b1;
            15'b00110101_0100_001: DATA = 1'b1;
            15'b00110101_0100_010: DATA = 1'b1;
            15'b00110101_0100_011: DATA = 1'b1;
            15'b00110101_0100_100: DATA = 1'b1;
            15'b00110101_0100_101: DATA = 1'b1;
            15'b00110101_0100_110: DATA = 1'b1;
            15'b00110101_0100_111: DATA = 1'b0;
            // 5 Row 5
            15'b00110101_0101_000: DATA = 1'b1;
            15'b00110101_0101_001: DATA = 1'b1;
            15'b00110101_0101_010: DATA = 1'b0;
            15'b00110101_0101_011: DATA = 1'b0;
            15'b00110101_0101_100: DATA = 1'b0;
            15'b00110101_0101_101: DATA = 1'b0;
            15'b00110101_0101_110: DATA = 1'b0;
            15'b00110101_0101_111: DATA = 1'b0;
            // 5 Row 6
            15'b00110101_0110_000: DATA = 1'b1;
            15'b00110101_0110_001: DATA = 1'b1;
            15'b00110101_0110_010: DATA = 1'b0;
            15'b00110101_0110_011: DATA = 1'b0;
            15'b00110101_0110_100: DATA = 1'b0;
            15'b00110101_0110_101: DATA = 1'b0;
            15'b00110101_0110_110: DATA = 1'b0;
            15'b00110101_0110_111: DATA = 1'b0;
            // 5 Row 7
            15'b00110101_0111_000: DATA = 1'b1;
            15'b00110101_0111_001: DATA = 1'b1;
            15'b00110101_0111_010: DATA = 1'b1;
            15'b00110101_0111_011: DATA = 1'b1;
            15'b00110101_0111_100: DATA = 1'b1;
            15'b00110101_0111_101: DATA = 1'b1;
            15'b00110101_0111_110: DATA = 1'b0;
            15'b00110101_0111_111: DATA = 1'b0;
            // 5 Row 8
            15'b00110101_1000_000: DATA = 1'b1;
            15'b00110101_1000_001: DATA = 1'b0;
            15'b00110101_1000_010: DATA = 1'b0;
            15'b00110101_1000_011: DATA = 1'b0;
            15'b00110101_1000_100: DATA = 1'b0;
            15'b00110101_1000_101: DATA = 1'b1;
            15'b00110101_1000_110: DATA = 1'b1;
            15'b00110101_1000_111: DATA = 1'b0;
            // 5 Row 9
            15'b00110101_1001_000: DATA = 1'b0;
            15'b00110101_1001_001: DATA = 1'b0;
            15'b00110101_1001_010: DATA = 1'b0;
            15'b00110101_1001_011: DATA = 1'b0;
            15'b00110101_1001_100: DATA = 1'b0;
            15'b00110101_1001_101: DATA = 1'b1;
            15'b00110101_1001_110: DATA = 1'b1;
            15'b00110101_1001_111: DATA = 1'b0;
            // 5 Row 10
            15'b00110101_1010_000: DATA = 1'b0;
            15'b00110101_1010_001: DATA = 1'b0;
            15'b00110101_1010_010: DATA = 1'b0;
            15'b00110101_1010_011: DATA = 1'b0;
            15'b00110101_1010_100: DATA = 1'b0;
            15'b00110101_1010_101: DATA = 1'b1;
            15'b00110101_1010_110: DATA = 1'b1;
            15'b00110101_1010_111: DATA = 1'b0;
            // 5 Row 11
            15'b00110101_1011_000: DATA = 1'b1;
            15'b00110101_1011_001: DATA = 1'b1;
            15'b00110101_1011_010: DATA = 1'b1;
            15'b00110101_1011_011: DATA = 1'b0;
            15'b00110101_1011_100: DATA = 1'b0;
            15'b00110101_1011_101: DATA = 1'b1;
            15'b00110101_1011_110: DATA = 1'b1;
            15'b00110101_1011_111: DATA = 1'b0;
            // 5 Row 12
            15'b00110101_1100_000: DATA = 1'b0;
            15'b00110101_1100_001: DATA = 1'b1;
            15'b00110101_1100_010: DATA = 1'b1;
            15'b00110101_1100_011: DATA = 1'b1;
            15'b00110101_1100_100: DATA = 1'b1;
            15'b00110101_1100_101: DATA = 1'b1;
            15'b00110101_1100_110: DATA = 1'b0;
            15'b00110101_1100_111: DATA = 1'b0;
            // 5 Row 13
            15'b00110101_1101_000: DATA = 1'b0;
            15'b00110101_1101_001: DATA = 1'b0;
            15'b00110101_1101_010: DATA = 1'b0;
            15'b00110101_1101_011: DATA = 1'b0;
            15'b00110101_1101_100: DATA = 1'b0;
            15'b00110101_1101_101: DATA = 1'b0;
            15'b00110101_1101_110: DATA = 1'b0;
            15'b00110101_1101_111: DATA = 1'b0;
            // 5 Row 14
            15'b00110101_1110_000: DATA = 1'b0;
            15'b00110101_1110_001: DATA = 1'b0;
            15'b00110101_1110_010: DATA = 1'b0;
            15'b00110101_1110_011: DATA = 1'b0;
            15'b00110101_1110_100: DATA = 1'b0;
            15'b00110101_1110_101: DATA = 1'b0;
            15'b00110101_1110_110: DATA = 1'b0;
            15'b00110101_1110_111: DATA = 1'b0;
            // 5 Row 15
            15'b00110101_1111_000: DATA = 1'b0;
            15'b00110101_1111_001: DATA = 1'b0;
            15'b00110101_1111_010: DATA = 1'b0;
            15'b00110101_1111_011: DATA = 1'b0;
            15'b00110101_1111_100: DATA = 1'b0;
            15'b00110101_1111_101: DATA = 1'b0;
            15'b00110101_1111_110: DATA = 1'b0;
            15'b00110101_1111_111: DATA = 1'b0;
            // 6 Row 0
            15'b00110110_0000_000: DATA = 1'b0;
            15'b00110110_0000_001: DATA = 1'b0;
            15'b00110110_0000_010: DATA = 1'b0;
            15'b00110110_0000_011: DATA = 1'b0;
            15'b00110110_0000_100: DATA = 1'b0;
            15'b00110110_0000_101: DATA = 1'b0;
            15'b00110110_0000_110: DATA = 1'b0;
            15'b00110110_0000_111: DATA = 1'b0;
            // 6 Row 1
            15'b00110110_0001_000: DATA = 1'b0;
            15'b00110110_0001_001: DATA = 1'b0;
            15'b00110110_0001_010: DATA = 1'b0;
            15'b00110110_0001_011: DATA = 1'b0;
            15'b00110110_0001_100: DATA = 1'b0;
            15'b00110110_0001_101: DATA = 1'b0;
            15'b00110110_0001_110: DATA = 1'b0;
            15'b00110110_0001_111: DATA = 1'b0;
            // 6 Row 2
            15'b00110110_0010_000: DATA = 1'b0;
            15'b00110110_0010_001: DATA = 1'b0;
            15'b00110110_0010_010: DATA = 1'b0;
            15'b00110110_0010_011: DATA = 1'b0;
            15'b00110110_0010_100: DATA = 1'b0;
            15'b00110110_0010_101: DATA = 1'b0;
            15'b00110110_0010_110: DATA = 1'b0;
            15'b00110110_0010_111: DATA = 1'b0;
            // 6 Row 3
            15'b00110110_0011_000: DATA = 1'b0;
            15'b00110110_0011_001: DATA = 1'b0;
            15'b00110110_0011_010: DATA = 1'b1;
            15'b00110110_0011_011: DATA = 1'b1;
            15'b00110110_0011_100: DATA = 1'b1;
            15'b00110110_0011_101: DATA = 1'b0;
            15'b00110110_0011_110: DATA = 1'b0;
            15'b00110110_0011_111: DATA = 1'b0;
            // 6 Row 4
            15'b00110110_0100_000: DATA = 1'b0;
            15'b00110110_0100_001: DATA = 1'b1;
            15'b00110110_0100_010: DATA = 1'b1;
            15'b00110110_0100_011: DATA = 1'b1;
            15'b00110110_0100_100: DATA = 1'b1;
            15'b00110110_0100_101: DATA = 1'b1;
            15'b00110110_0100_110: DATA = 1'b0;
            15'b00110110_0100_111: DATA = 1'b0;
            // 6 Row 5
            15'b00110110_0101_000: DATA = 1'b1;
            15'b00110110_0101_001: DATA = 1'b1;
            15'b00110110_0101_010: DATA = 1'b0;
            15'b00110110_0101_011: DATA = 1'b0;
            15'b00110110_0101_100: DATA = 1'b0;
            15'b00110110_0101_101: DATA = 1'b1;
            15'b00110110_0101_110: DATA = 1'b1;
            15'b00110110_0101_111: DATA = 1'b0;
            // 6 Row 6
            15'b00110110_0110_000: DATA = 1'b1;
            15'b00110110_0110_001: DATA = 1'b1;
            15'b00110110_0110_010: DATA = 1'b0;
            15'b00110110_0110_011: DATA = 1'b0;
            15'b00110110_0110_100: DATA = 1'b0;
            15'b00110110_0110_101: DATA = 1'b0;
            15'b00110110_0110_110: DATA = 1'b0;
            15'b00110110_0110_111: DATA = 1'b0;
            // 6 Row 7
            15'b00110110_0111_000: DATA = 1'b1;
            15'b00110110_0111_001: DATA = 1'b1;
            15'b00110110_0111_010: DATA = 1'b0;
            15'b00110110_0111_011: DATA = 1'b0;
            15'b00110110_0111_100: DATA = 1'b0;
            15'b00110110_0111_101: DATA = 1'b0;
            15'b00110110_0111_110: DATA = 1'b0;
            15'b00110110_0111_111: DATA = 1'b0;
            // 6 Row 8
            15'b00110110_1000_000: DATA = 1'b1;
            15'b00110110_1000_001: DATA = 1'b1;
            15'b00110110_1000_010: DATA = 1'b1;
            15'b00110110_1000_011: DATA = 1'b1;
            15'b00110110_1000_100: DATA = 1'b1;
            15'b00110110_1000_101: DATA = 1'b1;
            15'b00110110_1000_110: DATA = 1'b0;
            15'b00110110_1000_111: DATA = 1'b0;
            // 6 Row 9
            15'b00110110_1001_000: DATA = 1'b1;
            15'b00110110_1001_001: DATA = 1'b1;
            15'b00110110_1001_010: DATA = 1'b0;
            15'b00110110_1001_011: DATA = 1'b0;
            15'b00110110_1001_100: DATA = 1'b0;
            15'b00110110_1001_101: DATA = 1'b1;
            15'b00110110_1001_110: DATA = 1'b1;
            15'b00110110_1001_111: DATA = 1'b0;
            // 6 Row 10
            15'b00110110_1010_000: DATA = 1'b1;
            15'b00110110_1010_001: DATA = 1'b1;
            15'b00110110_1010_010: DATA = 1'b0;
            15'b00110110_1010_011: DATA = 1'b0;
            15'b00110110_1010_100: DATA = 1'b0;
            15'b00110110_1010_101: DATA = 1'b1;
            15'b00110110_1010_110: DATA = 1'b1;
            15'b00110110_1010_111: DATA = 1'b0;
            // 6 Row 11
            15'b00110110_1011_000: DATA = 1'b1;
            15'b00110110_1011_001: DATA = 1'b1;
            15'b00110110_1011_010: DATA = 1'b0;
            15'b00110110_1011_011: DATA = 1'b0;
            15'b00110110_1011_100: DATA = 1'b0;
            15'b00110110_1011_101: DATA = 1'b1;
            15'b00110110_1011_110: DATA = 1'b1;
            15'b00110110_1011_111: DATA = 1'b0;
            // 6 Row 12
            15'b00110110_1100_000: DATA = 1'b0;
            15'b00110110_1100_001: DATA = 1'b1;
            15'b00110110_1100_010: DATA = 1'b1;
            15'b00110110_1100_011: DATA = 1'b1;
            15'b00110110_1100_100: DATA = 1'b1;
            15'b00110110_1100_101: DATA = 1'b1;
            15'b00110110_1100_110: DATA = 1'b0;
            15'b00110110_1100_111: DATA = 1'b0;
            // 6 Row 13
            15'b00110110_1101_000: DATA = 1'b0;
            15'b00110110_1101_001: DATA = 1'b0;
            15'b00110110_1101_010: DATA = 1'b0;
            15'b00110110_1101_011: DATA = 1'b0;
            15'b00110110_1101_100: DATA = 1'b0;
            15'b00110110_1101_101: DATA = 1'b0;
            15'b00110110_1101_110: DATA = 1'b0;
            15'b00110110_1101_111: DATA = 1'b0;
            // 6 Row 14
            15'b00110110_1110_000: DATA = 1'b0;
            15'b00110110_1110_001: DATA = 1'b0;
            15'b00110110_1110_010: DATA = 1'b0;
            15'b00110110_1110_011: DATA = 1'b0;
            15'b00110110_1110_100: DATA = 1'b0;
            15'b00110110_1110_101: DATA = 1'b0;
            15'b00110110_1110_110: DATA = 1'b0;
            15'b00110110_1110_111: DATA = 1'b0;
            // 6 Row 15
            15'b00110110_1111_000: DATA = 1'b0;
            15'b00110110_1111_001: DATA = 1'b0;
            15'b00110110_1111_010: DATA = 1'b0;
            15'b00110110_1111_011: DATA = 1'b0;
            15'b00110110_1111_100: DATA = 1'b0;
            15'b00110110_1111_101: DATA = 1'b0;
            15'b00110110_1111_110: DATA = 1'b0;
            15'b00110110_1111_111: DATA = 1'b0;
            // 7 Row 0
            15'b00110111_0000_000: DATA = 1'b0;
            15'b00110111_0000_001: DATA = 1'b0;
            15'b00110111_0000_010: DATA = 1'b0;
            15'b00110111_0000_011: DATA = 1'b0;
            15'b00110111_0000_100: DATA = 1'b0;
            15'b00110111_0000_101: DATA = 1'b0;
            15'b00110111_0000_110: DATA = 1'b0;
            15'b00110111_0000_111: DATA = 1'b0;
            // 7 Row 1
            15'b00110111_0001_000: DATA = 1'b0;
            15'b00110111_0001_001: DATA = 1'b0;
            15'b00110111_0001_010: DATA = 1'b0;
            15'b00110111_0001_011: DATA = 1'b0;
            15'b00110111_0001_100: DATA = 1'b0;
            15'b00110111_0001_101: DATA = 1'b0;
            15'b00110111_0001_110: DATA = 1'b0;
            15'b00110111_0001_111: DATA = 1'b0;
            // 7 Row 2
            15'b00110111_0010_000: DATA = 1'b0;
            15'b00110111_0010_001: DATA = 1'b0;
            15'b00110111_0010_010: DATA = 1'b0;
            15'b00110111_0010_011: DATA = 1'b0;
            15'b00110111_0010_100: DATA = 1'b0;
            15'b00110111_0010_101: DATA = 1'b0;
            15'b00110111_0010_110: DATA = 1'b0;
            15'b00110111_0010_111: DATA = 1'b0;
            // 7 Row 3
            15'b00110111_0011_000: DATA = 1'b1;
            15'b00110111_0011_001: DATA = 1'b1;
            15'b00110111_0011_010: DATA = 1'b1;
            15'b00110111_0011_011: DATA = 1'b1;
            15'b00110111_0011_100: DATA = 1'b1;
            15'b00110111_0011_101: DATA = 1'b1;
            15'b00110111_0011_110: DATA = 1'b1;
            15'b00110111_0011_111: DATA = 1'b0;
            // 7 Row 4
            15'b00110111_0100_000: DATA = 1'b1;
            15'b00110111_0100_001: DATA = 1'b1;
            15'b00110111_0100_010: DATA = 1'b1;
            15'b00110111_0100_011: DATA = 1'b1;
            15'b00110111_0100_100: DATA = 1'b1;
            15'b00110111_0100_101: DATA = 1'b1;
            15'b00110111_0100_110: DATA = 1'b1;
            15'b00110111_0100_111: DATA = 1'b0;
            // 7 Row 5
            15'b00110111_0101_000: DATA = 1'b0;
            15'b00110111_0101_001: DATA = 1'b0;
            15'b00110111_0101_010: DATA = 1'b0;
            15'b00110111_0101_011: DATA = 1'b0;
            15'b00110111_0101_100: DATA = 1'b0;
            15'b00110111_0101_101: DATA = 1'b1;
            15'b00110111_0101_110: DATA = 1'b1;
            15'b00110111_0101_111: DATA = 1'b0;
            // 7 Row 6
            15'b00110111_0110_000: DATA = 1'b0;
            15'b00110111_0110_001: DATA = 1'b0;
            15'b00110111_0110_010: DATA = 1'b0;
            15'b00110111_0110_011: DATA = 1'b0;
            15'b00110111_0110_100: DATA = 1'b1;
            15'b00110111_0110_101: DATA = 1'b1;
            15'b00110111_0110_110: DATA = 1'b0;
            15'b00110111_0110_111: DATA = 1'b0;
            // 7 Row 7
            15'b00110111_0111_000: DATA = 1'b0;
            15'b00110111_0111_001: DATA = 1'b0;
            15'b00110111_0111_010: DATA = 1'b0;
            15'b00110111_0111_011: DATA = 1'b0;
            15'b00110111_0111_100: DATA = 1'b0;
            15'b00110111_0111_101: DATA = 1'b0;
            15'b00110111_0111_110: DATA = 1'b0;
            15'b00110111_0111_111: DATA = 1'b0;
            // 7 Row 8
            15'b00110111_1000_000: DATA = 1'b0;
            15'b00110111_1000_001: DATA = 1'b0;
            15'b00110111_1000_010: DATA = 1'b0;
            15'b00110111_1000_011: DATA = 1'b1;
            15'b00110111_1000_100: DATA = 1'b1;
            15'b00110111_1000_101: DATA = 1'b0;
            15'b00110111_1000_110: DATA = 1'b0;
            15'b00110111_1000_111: DATA = 1'b0;
            // 7 Row 9
            15'b00110111_1001_000: DATA = 1'b0;
            15'b00110111_1001_001: DATA = 1'b0;
            15'b00110111_1001_010: DATA = 1'b1;
            15'b00110111_1001_011: DATA = 1'b1;
            15'b00110111_1001_100: DATA = 1'b0;
            15'b00110111_1001_101: DATA = 1'b0;
            15'b00110111_1001_110: DATA = 1'b0;
            15'b00110111_1001_111: DATA = 1'b0;
            // 7 Row 10
            15'b00110111_1010_000: DATA = 1'b0;
            15'b00110111_1010_001: DATA = 1'b0;
            15'b00110111_1010_010: DATA = 1'b1;
            15'b00110111_1010_011: DATA = 1'b1;
            15'b00110111_1010_100: DATA = 1'b0;
            15'b00110111_1010_101: DATA = 1'b0;
            15'b00110111_1010_110: DATA = 1'b0;
            15'b00110111_1010_111: DATA = 1'b0;
            // 7 Row 11
            15'b00110111_1011_000: DATA = 1'b0;
            15'b00110111_1011_001: DATA = 1'b0;
            15'b00110111_1011_010: DATA = 1'b1;
            15'b00110111_1011_011: DATA = 1'b1;
            15'b00110111_1011_100: DATA = 1'b0;
            15'b00110111_1011_101: DATA = 1'b0;
            15'b00110111_1011_110: DATA = 1'b0;
            15'b00110111_1011_111: DATA = 1'b0;
            // 7 Row 12
            15'b00110111_1100_000: DATA = 1'b0;
            15'b00110111_1100_001: DATA = 1'b0;
            15'b00110111_1100_010: DATA = 1'b1;
            15'b00110111_1100_011: DATA = 1'b1;
            15'b00110111_1100_100: DATA = 1'b0;
            15'b00110111_1100_101: DATA = 1'b0;
            15'b00110111_1100_110: DATA = 1'b0;
            15'b00110111_1100_111: DATA = 1'b0;
            // 7 Row 13
            15'b00110111_1101_000: DATA = 1'b0;
            15'b00110111_1101_001: DATA = 1'b0;
            15'b00110111_1101_010: DATA = 1'b0;
            15'b00110111_1101_011: DATA = 1'b0;
            15'b00110111_1101_100: DATA = 1'b0;
            15'b00110111_1101_101: DATA = 1'b0;
            15'b00110111_1101_110: DATA = 1'b0;
            15'b00110111_1101_111: DATA = 1'b0;
            // 7 Row 14
            15'b00110111_1110_000: DATA = 1'b0;
            15'b00110111_1110_001: DATA = 1'b0;
            15'b00110111_1110_010: DATA = 1'b0;
            15'b00110111_1110_011: DATA = 1'b0;
            15'b00110111_1110_100: DATA = 1'b0;
            15'b00110111_1110_101: DATA = 1'b0;
            15'b00110111_1110_110: DATA = 1'b0;
            15'b00110111_1110_111: DATA = 1'b0;
            // 7 Row 15
            15'b00110111_1111_000: DATA = 1'b0;
            15'b00110111_1111_001: DATA = 1'b0;
            15'b00110111_1111_010: DATA = 1'b0;
            15'b00110111_1111_011: DATA = 1'b0;
            15'b00110111_1111_100: DATA = 1'b0;
            15'b00110111_1111_101: DATA = 1'b0;
            15'b00110111_1111_110: DATA = 1'b0;
            15'b00110111_1111_111: DATA = 1'b0;
            // 8 Row 0
            15'b00111000_0000_000: DATA = 1'b0;
            15'b00111000_0000_001: DATA = 1'b0;
            15'b00111000_0000_010: DATA = 1'b0;
            15'b00111000_0000_011: DATA = 1'b0;
            15'b00111000_0000_100: DATA = 1'b0;
            15'b00111000_0000_101: DATA = 1'b0;
            15'b00111000_0000_110: DATA = 1'b0;
            15'b00111000_0000_111: DATA = 1'b0;
            // 8 Row 1
            15'b00111000_0001_000: DATA = 1'b0;
            15'b00111000_0001_001: DATA = 1'b0;
            15'b00111000_0001_010: DATA = 1'b0;
            15'b00111000_0001_011: DATA = 1'b0;
            15'b00111000_0001_100: DATA = 1'b0;
            15'b00111000_0001_101: DATA = 1'b0;
            15'b00111000_0001_110: DATA = 1'b0;
            15'b00111000_0001_111: DATA = 1'b0;
            // 8 Row 2
            15'b00111000_0010_000: DATA = 1'b0;
            15'b00111000_0010_001: DATA = 1'b0;
            15'b00111000_0010_010: DATA = 1'b0;
            15'b00111000_0010_011: DATA = 1'b0;
            15'b00111000_0010_100: DATA = 1'b0;
            15'b00111000_0010_101: DATA = 1'b0;
            15'b00111000_0010_110: DATA = 1'b0;
            15'b00111000_0010_111: DATA = 1'b0;
            // 8 Row 3
            15'b00111000_0011_000: DATA = 1'b0;
            15'b00111000_0011_001: DATA = 1'b1;
            15'b00111000_0011_010: DATA = 1'b1;
            15'b00111000_0011_011: DATA = 1'b1;
            15'b00111000_0011_100: DATA = 1'b1;
            15'b00111000_0011_101: DATA = 1'b1;
            15'b00111000_0011_110: DATA = 1'b0;
            15'b00111000_0011_111: DATA = 1'b0;
            // 8 Row 4
            15'b00111000_0100_000: DATA = 1'b1;
            15'b00111000_0100_001: DATA = 1'b1;
            15'b00111000_0100_010: DATA = 1'b1;
            15'b00111000_0100_011: DATA = 1'b1;
            15'b00111000_0100_100: DATA = 1'b1;
            15'b00111000_0100_101: DATA = 1'b1;
            15'b00111000_0100_110: DATA = 1'b1;
            15'b00111000_0100_111: DATA = 1'b0;
            // 8 Row 5
            15'b00111000_0101_000: DATA = 1'b1;
            15'b00111000_0101_001: DATA = 1'b1;
            15'b00111000_0101_010: DATA = 1'b0;
            15'b00111000_0101_011: DATA = 1'b0;
            15'b00111000_0101_100: DATA = 1'b0;
            15'b00111000_0101_101: DATA = 1'b1;
            15'b00111000_0101_110: DATA = 1'b1;
            15'b00111000_0101_111: DATA = 1'b0;
            // 8 Row 6
            15'b00111000_0110_000: DATA = 1'b1;
            15'b00111000_0110_001: DATA = 1'b1;
            15'b00111000_0110_010: DATA = 1'b0;
            15'b00111000_0110_011: DATA = 1'b0;
            15'b00111000_0110_100: DATA = 1'b0;
            15'b00111000_0110_101: DATA = 1'b1;
            15'b00111000_0110_110: DATA = 1'b1;
            15'b00111000_0110_111: DATA = 1'b0;
            // 8 Row 7
            15'b00111000_0111_000: DATA = 1'b0;
            15'b00111000_0111_001: DATA = 1'b1;
            15'b00111000_0111_010: DATA = 1'b1;
            15'b00111000_0111_011: DATA = 1'b1;
            15'b00111000_0111_100: DATA = 1'b1;
            15'b00111000_0111_101: DATA = 1'b1;
            15'b00111000_0111_110: DATA = 1'b0;
            15'b00111000_0111_111: DATA = 1'b0;
            // 8 Row 8
            15'b00111000_1000_000: DATA = 1'b0;
            15'b00111000_1000_001: DATA = 1'b1;
            15'b00111000_1000_010: DATA = 1'b1;
            15'b00111000_1000_011: DATA = 1'b1;
            15'b00111000_1000_100: DATA = 1'b1;
            15'b00111000_1000_101: DATA = 1'b1;
            15'b00111000_1000_110: DATA = 1'b0;
            15'b00111000_1000_111: DATA = 1'b0;
            // 8 Row 9
            15'b00111000_1001_000: DATA = 1'b1;
            15'b00111000_1001_001: DATA = 1'b1;
            15'b00111000_1001_010: DATA = 1'b0;
            15'b00111000_1001_011: DATA = 1'b0;
            15'b00111000_1001_100: DATA = 1'b0;
            15'b00111000_1001_101: DATA = 1'b1;
            15'b00111000_1001_110: DATA = 1'b1;
            15'b00111000_1001_111: DATA = 1'b0;
            // 8 Row 10
            15'b00111000_1010_000: DATA = 1'b1;
            15'b00111000_1010_001: DATA = 1'b1;
            15'b00111000_1010_010: DATA = 1'b0;
            15'b00111000_1010_011: DATA = 1'b0;
            15'b00111000_1010_100: DATA = 1'b0;
            15'b00111000_1010_101: DATA = 1'b1;
            15'b00111000_1010_110: DATA = 1'b1;
            15'b00111000_1010_111: DATA = 1'b0;
            // 8 Row 11
            15'b00111000_1011_000: DATA = 1'b1;
            15'b00111000_1011_001: DATA = 1'b1;
            15'b00111000_1011_010: DATA = 1'b1;
            15'b00111000_1011_011: DATA = 1'b1;
            15'b00111000_1011_100: DATA = 1'b1;
            15'b00111000_1011_101: DATA = 1'b1;
            15'b00111000_1011_110: DATA = 1'b1;
            15'b00111000_1011_111: DATA = 1'b0;
            // 8 Row 12
            15'b00111000_1100_000: DATA = 1'b0;
            15'b00111000_1100_001: DATA = 1'b1;
            15'b00111000_1100_010: DATA = 1'b1;
            15'b00111000_1100_011: DATA = 1'b1;
            15'b00111000_1100_100: DATA = 1'b1;
            15'b00111000_1100_101: DATA = 1'b1;
            15'b00111000_1100_110: DATA = 1'b0;
            15'b00111000_1100_111: DATA = 1'b0;
            // 8 Row 13
            15'b00111000_1101_000: DATA = 1'b0;
            15'b00111000_1101_001: DATA = 1'b0;
            15'b00111000_1101_010: DATA = 1'b0;
            15'b00111000_1101_011: DATA = 1'b0;
            15'b00111000_1101_100: DATA = 1'b0;
            15'b00111000_1101_101: DATA = 1'b0;
            15'b00111000_1101_110: DATA = 1'b0;
            15'b00111000_1101_111: DATA = 1'b0;
            // 8 Row 14
            15'b00111000_1110_000: DATA = 1'b0;
            15'b00111000_1110_001: DATA = 1'b0;
            15'b00111000_1110_010: DATA = 1'b0;
            15'b00111000_1110_011: DATA = 1'b0;
            15'b00111000_1110_100: DATA = 1'b0;
            15'b00111000_1110_101: DATA = 1'b0;
            15'b00111000_1110_110: DATA = 1'b0;
            15'b00111000_1110_111: DATA = 1'b0;
            // 8 Row 15
            15'b00111000_1111_000: DATA = 1'b0;
            15'b00111000_1111_001: DATA = 1'b0;
            15'b00111000_1111_010: DATA = 1'b0;
            15'b00111000_1111_011: DATA = 1'b0;
            15'b00111000_1111_100: DATA = 1'b0;
            15'b00111000_1111_101: DATA = 1'b0;
            15'b00111000_1111_110: DATA = 1'b0;
            15'b00111000_1111_111: DATA = 1'b0;
            // 9 Row 0
            15'b00111001_0000_000: DATA = 1'b0;
            15'b00111001_0000_001: DATA = 1'b0;
            15'b00111001_0000_010: DATA = 1'b0;
            15'b00111001_0000_011: DATA = 1'b0;
            15'b00111001_0000_100: DATA = 1'b0;
            15'b00111001_0000_101: DATA = 1'b0;
            15'b00111001_0000_110: DATA = 1'b0;
            15'b00111001_0000_111: DATA = 1'b0;
            // 9 Row 1
            15'b00111001_0001_000: DATA = 1'b0;
            15'b00111001_0001_001: DATA = 1'b0;
            15'b00111001_0001_010: DATA = 1'b0;
            15'b00111001_0001_011: DATA = 1'b0;
            15'b00111001_0001_100: DATA = 1'b0;
            15'b00111001_0001_101: DATA = 1'b0;
            15'b00111001_0001_110: DATA = 1'b0;
            15'b00111001_0001_111: DATA = 1'b0;
            // 9 Row 2
            15'b00111001_0010_000: DATA = 1'b0;
            15'b00111001_0010_001: DATA = 1'b0;
            15'b00111001_0010_010: DATA = 1'b0;
            15'b00111001_0010_011: DATA = 1'b0;
            15'b00111001_0010_100: DATA = 1'b0;
            15'b00111001_0010_101: DATA = 1'b0;
            15'b00111001_0010_110: DATA = 1'b0;
            15'b00111001_0010_111: DATA = 1'b0;
            // 9 Row 3
            15'b00111001_0011_000: DATA = 1'b0;
            15'b00111001_0011_001: DATA = 1'b1;
            15'b00111001_0011_010: DATA = 1'b1;
            15'b00111001_0011_011: DATA = 1'b1;
            15'b00111001_0011_100: DATA = 1'b1;
            15'b00111001_0011_101: DATA = 1'b1;
            15'b00111001_0011_110: DATA = 1'b0;
            15'b00111001_0011_111: DATA = 1'b0;
            // 9 Row 4
            15'b00111001_0100_000: DATA = 1'b1;
            15'b00111001_0100_001: DATA = 1'b1;
            15'b00111001_0100_010: DATA = 1'b1;
            15'b00111001_0100_011: DATA = 1'b1;
            15'b00111001_0100_100: DATA = 1'b1;
            15'b00111001_0100_101: DATA = 1'b1;
            15'b00111001_0100_110: DATA = 1'b1;
            15'b00111001_0100_111: DATA = 1'b0;
            // 9 Row 5
            15'b00111001_0101_000: DATA = 1'b1;
            15'b00111001_0101_001: DATA = 1'b1;
            15'b00111001_0101_010: DATA = 1'b0;
            15'b00111001_0101_011: DATA = 1'b0;
            15'b00111001_0101_100: DATA = 1'b0;
            15'b00111001_0101_101: DATA = 1'b1;
            15'b00111001_0101_110: DATA = 1'b1;
            15'b00111001_0101_111: DATA = 1'b0;
            // 9 Row 6
            15'b00111001_0110_000: DATA = 1'b1;
            15'b00111001_0110_001: DATA = 1'b1;
            15'b00111001_0110_010: DATA = 1'b0;
            15'b00111001_0110_011: DATA = 1'b0;
            15'b00111001_0110_100: DATA = 1'b0;
            15'b00111001_0110_101: DATA = 1'b1;
            15'b00111001_0110_110: DATA = 1'b1;
            15'b00111001_0110_111: DATA = 1'b0;
            // 9 Row 7
            15'b00111001_0111_000: DATA = 1'b1;
            15'b00111001_0111_001: DATA = 1'b1;
            15'b00111001_0111_010: DATA = 1'b1;
            15'b00111001_0111_011: DATA = 1'b1;
            15'b00111001_0111_100: DATA = 1'b1;
            15'b00111001_0111_101: DATA = 1'b1;
            15'b00111001_0111_110: DATA = 1'b1;
            15'b00111001_0111_111: DATA = 1'b0;
            // 9 Row 8
            15'b00111001_1000_000: DATA = 1'b0;
            15'b00111001_1000_001: DATA = 1'b1;
            15'b00111001_1000_010: DATA = 1'b1;
            15'b00111001_1000_011: DATA = 1'b1;
            15'b00111001_1000_100: DATA = 1'b1;
            15'b00111001_1000_101: DATA = 1'b1;
            15'b00111001_1000_110: DATA = 1'b1;
            15'b00111001_1000_111: DATA = 1'b0;
            // 9 Row 9
            15'b00111001_1001_000: DATA = 1'b0;
            15'b00111001_1001_001: DATA = 1'b0;
            15'b00111001_1001_010: DATA = 1'b0;
            15'b00111001_1001_011: DATA = 1'b0;
            15'b00111001_1001_100: DATA = 1'b0;
            15'b00111001_1001_101: DATA = 1'b1;
            15'b00111001_1001_110: DATA = 1'b1;
            15'b00111001_1001_111: DATA = 1'b0;
            // 9 Row 10
            15'b00111001_1010_000: DATA = 1'b1;
            15'b00111001_1010_001: DATA = 1'b0;
            15'b00111001_1010_010: DATA = 1'b0;
            15'b00111001_1010_011: DATA = 1'b0;
            15'b00111001_1010_100: DATA = 1'b0;
            15'b00111001_1010_101: DATA = 1'b1;
            15'b00111001_1010_110: DATA = 1'b1;
            15'b00111001_1010_111: DATA = 1'b0;
            // < Row 0
            15'b00111100_0000_000: DATA = 1'b0;
            15'b00111100_0000_001: DATA = 1'b0;
            15'b00111100_0000_010: DATA = 1'b0;
            15'b00111100_0000_011: DATA = 1'b0;
            15'b00111100_0000_100: DATA = 1'b0;
            15'b00111100_0000_101: DATA = 1'b0;
            15'b00111100_0000_110: DATA = 1'b0;
            15'b00111100_0000_111: DATA = 1'b0;
            // < Row 1
            15'b00111100_0001_000: DATA = 1'b0;
            15'b00111100_0001_001: DATA = 1'b0;
            15'b00111100_0001_010: DATA = 1'b0;
            15'b00111100_0001_011: DATA = 1'b0;
            15'b00111100_0001_100: DATA = 1'b0;
            15'b00111100_0001_101: DATA = 1'b0;
            15'b00111100_0001_110: DATA = 1'b0;
            15'b00111100_0001_111: DATA = 1'b0;
            // < Row 2
            15'b00111100_0010_000: DATA = 1'b0;
            15'b00111100_0010_001: DATA = 1'b0;
            15'b00111100_0010_010: DATA = 1'b0;
            15'b00111100_0010_011: DATA = 1'b0;
            15'b00111100_0010_100: DATA = 1'b0;
            15'b00111100_0010_101: DATA = 1'b0;
            15'b00111100_0010_110: DATA = 1'b0;
            15'b00111100_0010_111: DATA = 1'b0;
            // < Row 3
            15'b00111100_0011_000: DATA = 1'b0;
            15'b00111100_0011_001: DATA = 1'b0;
            15'b00111100_0011_010: DATA = 1'b0;
            15'b00111100_0011_011: DATA = 1'b0;
            15'b00111100_0011_100: DATA = 1'b0;
            15'b00111100_0011_101: DATA = 1'b0;
            15'b00111100_0011_110: DATA = 1'b0;
            15'b00111100_0011_111: DATA = 1'b0;
            // < Row 4
            15'b00111100_0100_000: DATA = 1'b0;
            15'b00111100_0100_001: DATA = 1'b0;
            15'b00111100_0100_010: DATA = 1'b0;
            15'b00111100_0100_011: DATA = 1'b0;
            15'b00111100_0100_100: DATA = 1'b1;
            15'b00111100_0100_101: DATA = 1'b1;
            15'b00111100_0100_110: DATA = 1'b0;
            15'b00111100_0100_111: DATA = 1'b0;
            // < Row 5
            15'b00111100_0101_000: DATA = 1'b0;
            15'b00111100_0101_001: DATA = 1'b0;
            15'b00111100_0101_010: DATA = 1'b0;
            15'b00111100_0101_011: DATA = 1'b1;
            15'b00111100_0101_100: DATA = 1'b1;
            15'b00111100_0101_101: DATA = 1'b0;
            15'b00111100_0101_110: DATA = 1'b0;
            15'b00111100_0101_111: DATA = 1'b0;
            // < Row 6
            15'b00111100_0110_000: DATA = 1'b0;
            15'b00111100_0110_001: DATA = 1'b0;
            15'b00111100_0110_010: DATA = 1'b1;
            15'b00111100_0110_011: DATA = 1'b1;
            15'b00111100_0110_100: DATA = 1'b0;
            15'b00111100_0110_101: DATA = 1'b0;
            15'b00111100_0110_110: DATA = 1'b0;
            15'b00111100_0110_111: DATA = 1'b0;
            // < Row 7
            15'b00111100_0111_000: DATA = 1'b0;
            15'b00111100_0111_001: DATA = 1'b1;
            15'b00111100_0111_010: DATA = 1'b1;
            15'b00111100_0111_011: DATA = 1'b0;
            15'b00111100_0111_100: DATA = 1'b0;
            15'b00111100_0111_101: DATA = 1'b0;
            15'b00111100_0111_110: DATA = 1'b0;
            15'b00111100_0111_111: DATA = 1'b0;
            // < Row 8
            15'b00111100_1000_000: DATA = 1'b0;
            15'b00111100_1000_001: DATA = 1'b1;
            15'b00111100_1000_010: DATA = 1'b1;
            15'b00111100_1000_011: DATA = 1'b0;
            15'b00111100_1000_100: DATA = 1'b0;
            15'b00111100_1000_101: DATA = 1'b0;
            15'b00111100_1000_110: DATA = 1'b0;
            15'b00111100_1000_111: DATA = 1'b0;
            // < Row 9
            15'b00111100_1001_000: DATA = 1'b0;
            15'b00111100_1001_001: DATA = 1'b0;
            15'b00111100_1001_010: DATA = 1'b1;
            15'b00111100_1001_011: DATA = 1'b1;
            15'b00111100_1001_100: DATA = 1'b0;
            15'b00111100_1001_101: DATA = 1'b0;
            15'b00111100_1001_110: DATA = 1'b0;
            15'b00111100_1001_111: DATA = 1'b0;
            // < Row 10
            15'b00111100_1010_000: DATA = 1'b0;
            15'b00111100_1010_001: DATA = 1'b0;
            15'b00111100_1010_010: DATA = 1'b0;
            15'b00111100_1010_011: DATA = 1'b1;
            15'b00111100_1010_100: DATA = 1'b1;
            15'b00111100_1010_101: DATA = 1'b0;
            15'b00111100_1010_110: DATA = 1'b0;
            15'b00111100_1010_111: DATA = 1'b0;
            // < Row 11
            15'b00111100_1011_000: DATA = 1'b0;
            15'b00111100_1011_001: DATA = 1'b0;
            15'b00111100_1011_010: DATA = 1'b0;
            15'b00111100_1011_011: DATA = 1'b0;
            15'b00111100_1011_100: DATA = 1'b1;
            15'b00111100_1011_101: DATA = 1'b1;
            15'b00111100_1011_110: DATA = 1'b0;
            15'b00111100_1011_111: DATA = 1'b0;
            // < Row 12
            15'b00111100_1100_000: DATA = 1'b0;
            15'b00111100_1100_001: DATA = 1'b0;
            15'b00111100_1100_010: DATA = 1'b0;
            15'b00111100_1100_011: DATA = 1'b0;
            15'b00111100_1100_100: DATA = 1'b0;
            15'b00111100_1100_101: DATA = 1'b0;
            15'b00111100_1100_110: DATA = 1'b0;
            15'b00111100_1100_111: DATA = 1'b0;
            // < Row 13
            15'b00111100_1101_000: DATA = 1'b0;
            15'b00111100_1101_001: DATA = 1'b0;
            15'b00111100_1101_010: DATA = 1'b0;
            15'b00111100_1101_011: DATA = 1'b0;
            15'b00111100_1101_100: DATA = 1'b0;
            15'b00111100_1101_101: DATA = 1'b0;
            15'b00111100_1101_110: DATA = 1'b0;
            15'b00111100_1101_111: DATA = 1'b0;
            // < Row 14
            15'b00111100_1110_000: DATA = 1'b0;
            15'b00111100_1110_001: DATA = 1'b0;
            15'b00111100_1110_010: DATA = 1'b0;
            15'b00111100_1110_011: DATA = 1'b0;
            15'b00111100_1110_100: DATA = 1'b0;
            15'b00111100_1110_101: DATA = 1'b0;
            15'b00111100_1110_110: DATA = 1'b0;
            15'b00111100_1110_111: DATA = 1'b0;
            // < Row 15
            15'b00111100_1111_000: DATA = 1'b0;
            15'b00111100_1111_001: DATA = 1'b0;
            15'b00111100_1111_010: DATA = 1'b0;
            15'b00111100_1111_011: DATA = 1'b0;
            15'b00111100_1111_100: DATA = 1'b0;
            15'b00111100_1111_101: DATA = 1'b0;
            15'b00111100_1111_110: DATA = 1'b0;
            15'b00111100_1111_111: DATA = 1'b0;
            // 9 Row 11
            15'b00111001_1011_000: DATA = 1'b1;
            15'b00111001_1011_001: DATA = 1'b1;
            15'b00111001_1011_010: DATA = 1'b0;
            15'b00111001_1011_011: DATA = 1'b0;
            15'b00111001_1011_100: DATA = 1'b0;
            15'b00111001_1011_101: DATA = 1'b1;
            15'b00111001_1011_110: DATA = 1'b1;
            15'b00111001_1011_111: DATA = 1'b0;
            // 9 Row 12
            15'b00111001_1100_000: DATA = 1'b0;
            15'b00111001_1100_001: DATA = 1'b1;
            15'b00111001_1100_010: DATA = 1'b1;
            15'b00111001_1100_011: DATA = 1'b1;
            15'b00111001_1100_100: DATA = 1'b1;
            15'b00111001_1100_101: DATA = 1'b1;
            15'b00111001_1100_110: DATA = 1'b0;
            15'b00111001_1100_111: DATA = 1'b0;
            // 9 Row 13
            15'b00111001_1101_000: DATA = 1'b0;
            15'b00111001_1101_001: DATA = 1'b0;
            15'b00111001_1101_010: DATA = 1'b0;
            15'b00111001_1101_011: DATA = 1'b0;
            15'b00111001_1101_100: DATA = 1'b0;
            15'b00111001_1101_101: DATA = 1'b0;
            15'b00111001_1101_110: DATA = 1'b0;
            15'b00111001_1101_111: DATA = 1'b0;
            // 9 Row 14
            15'b00111001_1110_000: DATA = 1'b0;
            15'b00111001_1110_001: DATA = 1'b0;
            15'b00111001_1110_010: DATA = 1'b0;
            15'b00111001_1110_011: DATA = 1'b0;
            15'b00111001_1110_100: DATA = 1'b0;
            15'b00111001_1110_101: DATA = 1'b0;
            15'b00111001_1110_110: DATA = 1'b0;
            15'b00111001_1110_111: DATA = 1'b0;
            // 9 Row 15
            15'b00111001_1111_000: DATA = 1'b0;
            15'b00111001_1111_001: DATA = 1'b0;
            15'b00111001_1111_010: DATA = 1'b0;
            15'b00111001_1111_011: DATA = 1'b0;
            15'b00111001_1111_100: DATA = 1'b0;
            15'b00111001_1111_101: DATA = 1'b0;
            15'b00111001_1111_110: DATA = 1'b0;
            15'b00111001_1111_111: DATA = 1'b0;
            // A Row 0
            15'b01000001_0000_000: DATA = 1'b0;
            15'b01000001_0000_001: DATA = 1'b0;
            15'b01000001_0000_010: DATA = 1'b0;
            15'b01000001_0000_011: DATA = 1'b0;
            15'b01000001_0000_100: DATA = 1'b0;
            15'b01000001_0000_101: DATA = 1'b0;
            15'b01000001_0000_110: DATA = 1'b0;
            15'b01000001_0000_111: DATA = 1'b0;
            // A Row 1
            15'b01000001_0001_000: DATA = 1'b0;
            15'b01000001_0001_001: DATA = 1'b0;
            15'b01000001_0001_010: DATA = 1'b0;
            15'b01000001_0001_011: DATA = 1'b0;
            15'b01000001_0001_100: DATA = 1'b0;
            15'b01000001_0001_101: DATA = 1'b0;
            15'b01000001_0001_110: DATA = 1'b0;
            15'b01000001_0001_111: DATA = 1'b0;
            // A Row 2
            15'b01000001_0010_000: DATA = 1'b0;
            15'b01000001_0010_001: DATA = 1'b0;
            15'b01000001_0010_010: DATA = 1'b0;
            15'b01000001_0010_011: DATA = 1'b0;
            15'b01000001_0010_100: DATA = 1'b0;
            15'b01000001_0010_101: DATA = 1'b0;
            15'b01000001_0010_110: DATA = 1'b0;
            15'b01000001_0010_111: DATA = 1'b0;
            // A Row 3
            15'b01000001_0011_000: DATA = 1'b0;
            15'b01000001_0011_001: DATA = 1'b0;
            15'b01000001_0011_010: DATA = 1'b0;
            15'b01000001_0011_011: DATA = 1'b1;
            15'b01000001_0011_100: DATA = 1'b0;
            15'b01000001_0011_101: DATA = 1'b0;
            15'b01000001_0011_110: DATA = 1'b0;
            15'b01000001_0011_111: DATA = 1'b0;
            // A Row 4
            15'b01000001_0100_000: DATA = 1'b0;
            15'b01000001_0100_001: DATA = 1'b0;
            15'b01000001_0100_010: DATA = 1'b1;
            15'b01000001_0100_011: DATA = 1'b1;
            15'b01000001_0100_100: DATA = 1'b1;
            15'b01000001_0100_101: DATA = 1'b0;
            15'b01000001_0100_110: DATA = 1'b0;
            15'b01000001_0100_111: DATA = 1'b0;
            // A Row 5
            15'b01000001_0101_000: DATA = 1'b0;
            15'b01000001_0101_001: DATA = 1'b1;
            15'b01000001_0101_010: DATA = 1'b1;
            15'b01000001_0101_011: DATA = 1'b0;
            15'b01000001_0101_100: DATA = 1'b1;
            15'b01000001_0101_101: DATA = 1'b1;
            15'b01000001_0101_110: DATA = 1'b0;
            15'b01000001_0101_111: DATA = 1'b0;
            // A Row 6
            15'b01000001_0110_000: DATA = 1'b1;
            15'b01000001_0110_001: DATA = 1'b1;
            15'b01000001_0110_010: DATA = 1'b0;
            15'b01000001_0110_011: DATA = 1'b0;
            15'b01000001_0110_100: DATA = 1'b0;
            15'b01000001_0110_101: DATA = 1'b1;
            15'b01000001_0110_110: DATA = 1'b1;
            15'b01000001_0110_111: DATA = 1'b0;
            // A Row 7
            15'b01000001_0111_000: DATA = 1'b1;
            15'b01000001_0111_001: DATA = 1'b1;
            15'b01000001_0111_010: DATA = 1'b0;
            15'b01000001_0111_011: DATA = 1'b0;
            15'b01000001_0111_100: DATA = 1'b0;
            15'b01000001_0111_101: DATA = 1'b1;
            15'b01000001_0111_110: DATA = 1'b1;
            15'b01000001_0111_111: DATA = 1'b0;
            // A Row 8
            15'b01000001_1000_000: DATA = 1'b1;
            15'b01000001_1000_001: DATA = 1'b1;
            15'b01000001_1000_010: DATA = 1'b1;
            15'b01000001_1000_011: DATA = 1'b1;
            15'b01000001_1000_100: DATA = 1'b1;
            15'b01000001_1000_101: DATA = 1'b1;
            15'b01000001_1000_110: DATA = 1'b1;
            15'b01000001_1000_111: DATA = 1'b0;
            // A Row 9
            15'b01000001_1001_000: DATA = 1'b1;
            15'b01000001_1001_001: DATA = 1'b1;
            15'b01000001_1001_010: DATA = 1'b0;
            15'b01000001_1001_011: DATA = 1'b0;
            15'b01000001_1001_100: DATA = 1'b0;
            15'b01000001_1001_101: DATA = 1'b1;
            15'b01000001_1001_110: DATA = 1'b1;
            15'b01000001_1001_111: DATA = 1'b0;
            // A Row 10
            15'b01000001_1010_000: DATA = 1'b1;
            15'b01000001_1010_001: DATA = 1'b1;
            15'b01000001_1010_010: DATA = 1'b0;
            15'b01000001_1010_011: DATA = 1'b0;
            15'b01000001_1010_100: DATA = 1'b0;
            15'b01000001_1010_101: DATA = 1'b1;
            15'b01000001_1010_110: DATA = 1'b1;
            15'b01000001_1010_111: DATA = 1'b0;
            // A Row 11
            15'b01000001_1011_000: DATA = 1'b1;
            15'b01000001_1011_001: DATA = 1'b1;
            15'b01000001_1011_010: DATA = 1'b0;
            15'b01000001_1011_011: DATA = 1'b0;
            15'b01000001_1011_100: DATA = 1'b0;
            15'b01000001_1011_101: DATA = 1'b1;
            15'b01000001_1011_110: DATA = 1'b1;
            15'b01000001_1011_111: DATA = 1'b0;
            // A Row 12
            15'b01000001_1100_000: DATA = 1'b1;
            15'b01000001_1100_001: DATA = 1'b1;
            15'b01000001_1100_010: DATA = 1'b0;
            15'b01000001_1100_011: DATA = 1'b0;
            15'b01000001_1100_100: DATA = 1'b0;
            15'b01000001_1100_101: DATA = 1'b1;
            15'b01000001_1100_110: DATA = 1'b1;
            15'b01000001_1100_111: DATA = 1'b0;
            // A Row 13
            15'b01000001_1101_000: DATA = 1'b0;
            15'b01000001_1101_001: DATA = 1'b0;
            15'b01000001_1101_010: DATA = 1'b0;
            15'b01000001_1101_011: DATA = 1'b0;
            15'b01000001_1101_100: DATA = 1'b0;
            15'b01000001_1101_101: DATA = 1'b0;
            15'b01000001_1101_110: DATA = 1'b0;
            15'b01000001_1101_111: DATA = 1'b0;
            // A Row 14
            15'b01000001_1110_000: DATA = 1'b0;
            15'b01000001_1110_001: DATA = 1'b0;
            15'b01000001_1110_010: DATA = 1'b0;
            15'b01000001_1110_011: DATA = 1'b0;
            15'b01000001_1110_100: DATA = 1'b0;
            15'b01000001_1110_101: DATA = 1'b0;
            15'b01000001_1110_110: DATA = 1'b0;
            15'b01000001_1110_111: DATA = 1'b0;
            // A Row 15
            15'b01000001_1111_000: DATA = 1'b0;
            15'b01000001_1111_001: DATA = 1'b0;
            15'b01000001_1111_010: DATA = 1'b0;
            15'b01000001_1111_011: DATA = 1'b0;
            15'b01000001_1111_100: DATA = 1'b0;
            15'b01000001_1111_101: DATA = 1'b0;
            15'b01000001_1111_110: DATA = 1'b0;
            15'b01000001_1111_111: DATA = 1'b0;
            // B Row 0
            15'b01000010_0000_000: DATA = 1'b0;
            15'b01000010_0000_001: DATA = 1'b0;
            15'b01000010_0000_010: DATA = 1'b0;
            15'b01000010_0000_011: DATA = 1'b0;
            15'b01000010_0000_100: DATA = 1'b0;
            15'b01000010_0000_101: DATA = 1'b0;
            15'b01000010_0000_110: DATA = 1'b0;
            15'b01000010_0000_111: DATA = 1'b0;
            // B Row 1
            15'b01000010_0001_000: DATA = 1'b0;
            15'b01000010_0001_001: DATA = 1'b0;
            15'b01000010_0001_010: DATA = 1'b0;
            15'b01000010_0001_011: DATA = 1'b0;
            15'b01000010_0001_100: DATA = 1'b0;
            15'b01000010_0001_101: DATA = 1'b0;
            15'b01000010_0001_110: DATA = 1'b0;
            15'b01000010_0001_111: DATA = 1'b0;
            // B Row 2
            15'b01000010_0010_000: DATA = 1'b0;
            15'b01000010_0010_001: DATA = 1'b0;
            15'b01000010_0010_010: DATA = 1'b0;
            15'b01000010_0010_011: DATA = 1'b0;
            15'b01000010_0010_100: DATA = 1'b0;
            15'b01000010_0010_101: DATA = 1'b0;
            15'b01000010_0010_110: DATA = 1'b0;
            15'b01000010_0010_111: DATA = 1'b0;
            // B Row 3
            15'b01000010_0011_000: DATA = 1'b1;
            15'b01000010_0011_001: DATA = 1'b1;
            15'b01000010_0011_010: DATA = 1'b1;
            15'b01000010_0011_011: DATA = 1'b1;
            15'b01000010_0011_100: DATA = 1'b1;
            15'b01000010_0011_101: DATA = 1'b0;
            15'b01000010_0011_110: DATA = 1'b0;
            15'b01000010_0011_111: DATA = 1'b0;
            // B Row 4
            15'b01000010_0100_000: DATA = 1'b1;
            15'b01000010_0100_001: DATA = 1'b1;
            15'b01000010_0100_010: DATA = 1'b0;
            15'b01000010_0100_011: DATA = 1'b0;
            15'b01000010_0100_100: DATA = 1'b1;
            15'b01000010_0100_101: DATA = 1'b1;
            15'b01000010_0100_110: DATA = 1'b0;
            15'b01000010_0100_111: DATA = 1'b0;
            // B Row 5
            15'b01000010_0101_000: DATA = 1'b1;
            15'b01000010_0101_001: DATA = 1'b1;
            15'b01000010_0101_010: DATA = 1'b0;
            15'b01000010_0101_011: DATA = 1'b0;
            15'b01000010_0101_100: DATA = 1'b0;
            15'b01000010_0101_101: DATA = 1'b1;
            15'b01000010_0101_110: DATA = 1'b0;
            15'b01000010_0101_111: DATA = 1'b0;
            // B Row 6
            15'b01000010_0110_000: DATA = 1'b1;
            15'b01000010_0110_001: DATA = 1'b1;
            15'b01000010_0110_010: DATA = 1'b0;
            15'b01000010_0110_011: DATA = 1'b0;
            15'b01000010_0110_100: DATA = 1'b1;
            15'b01000010_0110_101: DATA = 1'b1;
            15'b01000010_0110_110: DATA = 1'b0;
            15'b01000010_0110_111: DATA = 1'b0;
            // B Row 7
            15'b01000010_0111_000: DATA = 1'b1;
            15'b01000010_0111_001: DATA = 1'b1;
            15'b01000010_0111_010: DATA = 1'b1;
            15'b01000010_0111_011: DATA = 1'b1;
            15'b01000010_0111_100: DATA = 1'b1;
            15'b01000010_0111_101: DATA = 1'b0;
            15'b01000010_0111_110: DATA = 1'b0;
            15'b01000010_0111_111: DATA = 1'b0;
            // B Row 8
            15'b01000010_1000_000: DATA = 1'b1;
            15'b01000010_1000_001: DATA = 1'b1;
            15'b01000010_1000_010: DATA = 1'b0;
            15'b01000010_1000_011: DATA = 1'b0;
            15'b01000010_1000_100: DATA = 1'b1;
            15'b01000010_1000_101: DATA = 1'b1;
            15'b01000010_1000_110: DATA = 1'b0;
            15'b01000010_1000_111: DATA = 1'b0;
            // B Row 9
            15'b01000010_1001_000: DATA = 1'b1;
            15'b01000010_1001_001: DATA = 1'b1;
            15'b01000010_1001_010: DATA = 1'b0;
            15'b01000010_1001_011: DATA = 1'b0;
            15'b01000010_1001_100: DATA = 1'b0;
            15'b01000010_1001_101: DATA = 1'b1;
            15'b01000010_1001_110: DATA = 1'b1;
            15'b01000010_1001_111: DATA = 1'b0;
            // B Row 10
            15'b01000010_1010_000: DATA = 1'b1;
            15'b01000010_1010_001: DATA = 1'b1;
            15'b01000010_1010_010: DATA = 1'b0;
            15'b01000010_1010_011: DATA = 1'b0;
            15'b01000010_1010_100: DATA = 1'b0;
            15'b01000010_1010_101: DATA = 1'b1;
            15'b01000010_1010_110: DATA = 1'b1;
            15'b01000010_1010_111: DATA = 1'b0;
            // B Row 11
            15'b01000010_1011_000: DATA = 1'b1;
            15'b01000010_1011_001: DATA = 1'b1;
            15'b01000010_1011_010: DATA = 1'b0;
            15'b01000010_1011_011: DATA = 1'b0;
            15'b01000010_1011_100: DATA = 1'b1;
            15'b01000010_1011_101: DATA = 1'b1;
            15'b01000010_1011_110: DATA = 1'b0;
            15'b01000010_1011_111: DATA = 1'b0;
            // B Row 12
            15'b01000010_1100_000: DATA = 1'b1;
            15'b01000010_1100_001: DATA = 1'b1;
            15'b01000010_1100_010: DATA = 1'b1;
            15'b01000010_1100_011: DATA = 1'b1;
            15'b01000010_1100_100: DATA = 1'b1;
            15'b01000010_1100_101: DATA = 1'b0;
            15'b01000010_1100_110: DATA = 1'b0;
            15'b01000010_1100_111: DATA = 1'b0;
            // B Row 13
            15'b01000010_1101_000: DATA = 1'b0;
            15'b01000010_1101_001: DATA = 1'b0;
            15'b01000010_1101_010: DATA = 1'b0;
            15'b01000010_1101_011: DATA = 1'b0;
            15'b01000010_1101_100: DATA = 1'b0;
            15'b01000010_1101_101: DATA = 1'b0;
            15'b01000010_1101_110: DATA = 1'b0;
            15'b01000010_1101_111: DATA = 1'b0;
            // B Row 14
            15'b01000010_1110_000: DATA = 1'b0;
            15'b01000010_1110_001: DATA = 1'b0;
            15'b01000010_1110_010: DATA = 1'b0;
            15'b01000010_1110_011: DATA = 1'b0;
            15'b01000010_1110_100: DATA = 1'b0;
            15'b01000010_1110_101: DATA = 1'b0;
            15'b01000010_1110_110: DATA = 1'b0;
            15'b01000010_1110_111: DATA = 1'b0;
            // B Row 15
            15'b01000010_1111_000: DATA = 1'b0;
            15'b01000010_1111_001: DATA = 1'b0;
            15'b01000010_1111_010: DATA = 1'b0;
            15'b01000010_1111_011: DATA = 1'b0;
            15'b01000010_1111_100: DATA = 1'b0;
            15'b01000010_1111_101: DATA = 1'b0;
            15'b01000010_1111_110: DATA = 1'b0;
            15'b01000010_1111_111: DATA = 1'b0;
            // C Row 0
            15'b01000011_0000_000: DATA = 1'b0;
            15'b01000011_0000_001: DATA = 1'b0;
            15'b01000011_0000_010: DATA = 1'b0;
            15'b01000011_0000_011: DATA = 1'b0;
            15'b01000011_0000_100: DATA = 1'b0;
            15'b01000011_0000_101: DATA = 1'b0;
            15'b01000011_0000_110: DATA = 1'b0;
            15'b01000011_0000_111: DATA = 1'b0;
            // C Row 1
            15'b01000011_0001_000: DATA = 1'b0;
            15'b01000011_0001_001: DATA = 1'b0;
            15'b01000011_0001_010: DATA = 1'b0;
            15'b01000011_0001_011: DATA = 1'b0;
            15'b01000011_0001_100: DATA = 1'b0;
            15'b01000011_0001_101: DATA = 1'b0;
            15'b01000011_0001_110: DATA = 1'b0;
            15'b01000011_0001_111: DATA = 1'b0;
            // C Row 2
            15'b01000011_0010_000: DATA = 1'b0;
            15'b01000011_0010_001: DATA = 1'b0;
            15'b01000011_0010_010: DATA = 1'b0;
            15'b01000011_0010_011: DATA = 1'b0;
            15'b01000011_0010_100: DATA = 1'b0;
            15'b01000011_0010_101: DATA = 1'b0;
            15'b01000011_0010_110: DATA = 1'b0;
            15'b01000011_0010_111: DATA = 1'b0;
            // C Row 3
            15'b01000011_0011_000: DATA = 1'b0;
            15'b01000011_0011_001: DATA = 1'b0;
            15'b01000011_0011_010: DATA = 1'b1;
            15'b01000011_0011_011: DATA = 1'b1;
            15'b01000011_0011_100: DATA = 1'b1;
            15'b01000011_0011_101: DATA = 1'b0;
            15'b01000011_0011_110: DATA = 1'b0;
            15'b01000011_0011_111: DATA = 1'b0;
            // C Row 4
            15'b01000011_0100_000: DATA = 1'b0;
            15'b01000011_0100_001: DATA = 1'b1;
            15'b01000011_0100_010: DATA = 1'b1;
            15'b01000011_0100_011: DATA = 1'b1;
            15'b01000011_0100_100: DATA = 1'b1;
            15'b01000011_0100_101: DATA = 1'b1;
            15'b01000011_0100_110: DATA = 1'b0;
            15'b01000011_0100_111: DATA = 1'b0;
            // C Row 5
            15'b01000011_0101_000: DATA = 1'b1;
            15'b01000011_0101_001: DATA = 1'b1;
            15'b01000011_0101_010: DATA = 1'b0;
            15'b01000011_0101_011: DATA = 1'b0;
            15'b01000011_0101_100: DATA = 1'b0;
            15'b01000011_0101_101: DATA = 1'b1;
            15'b01000011_0101_110: DATA = 1'b1;
            15'b01000011_0101_111: DATA = 1'b0;
            // C Row 6
            15'b01000011_0110_000: DATA = 1'b1;
            15'b01000011_0110_001: DATA = 1'b1;
            15'b01000011_0110_010: DATA = 1'b0;
            15'b01000011_0110_011: DATA = 1'b0;
            15'b01000011_0110_100: DATA = 1'b0;
            15'b01000011_0110_101: DATA = 1'b0;
            15'b01000011_0110_110: DATA = 1'b0;
            15'b01000011_0110_111: DATA = 1'b0;
            // C Row 7
            15'b01000011_0111_000: DATA = 1'b1;
            15'b01000011_0111_001: DATA = 1'b1;
            15'b01000011_0111_010: DATA = 1'b0;
            15'b01000011_0111_011: DATA = 1'b0;
            15'b01000011_0111_100: DATA = 1'b0;
            15'b01000011_0111_101: DATA = 1'b0;
            15'b01000011_0111_110: DATA = 1'b0;
            15'b01000011_0111_111: DATA = 1'b0;
            // C Row 8
            15'b01000011_1000_000: DATA = 1'b1;
            15'b01000011_1000_001: DATA = 1'b1;
            15'b01000011_1000_010: DATA = 1'b0;
            15'b01000011_1000_011: DATA = 1'b0;
            15'b01000011_1000_100: DATA = 1'b0;
            15'b01000011_1000_101: DATA = 1'b0;
            15'b01000011_1000_110: DATA = 1'b0;
            15'b01000011_1000_111: DATA = 1'b0;
            // C Row 9
            15'b01000011_1001_000: DATA = 1'b1;
            15'b01000011_1001_001: DATA = 1'b1;
            15'b01000011_1001_010: DATA = 1'b0;
            15'b01000011_1001_011: DATA = 1'b0;
            15'b01000011_1001_100: DATA = 1'b0;
            15'b01000011_1001_101: DATA = 1'b0;
            15'b01000011_1001_110: DATA = 1'b0;
            15'b01000011_1001_111: DATA = 1'b0;
            // C Row 10
            15'b01000011_1010_000: DATA = 1'b1;
            15'b01000011_1010_001: DATA = 1'b1;
            15'b01000011_1010_010: DATA = 1'b0;
            15'b01000011_1010_011: DATA = 1'b0;
            15'b01000011_1010_100: DATA = 1'b0;
            15'b01000011_1010_101: DATA = 1'b1;
            15'b01000011_1010_110: DATA = 1'b1;
            15'b01000011_1010_111: DATA = 1'b0;
            // C Row 11
            15'b01000011_1011_000: DATA = 1'b0;
            15'b01000011_1011_001: DATA = 1'b1;
            15'b01000011_1011_010: DATA = 1'b1;
            15'b01000011_1011_011: DATA = 1'b1;
            15'b01000011_1011_100: DATA = 1'b1;
            15'b01000011_1011_101: DATA = 1'b1;
            15'b01000011_1011_110: DATA = 1'b0;
            15'b01000011_1011_111: DATA = 1'b0;
            // C Row 12
            15'b01000011_1100_000: DATA = 1'b0;
            15'b01000011_1100_001: DATA = 1'b0;
            15'b01000011_1100_010: DATA = 1'b1;
            15'b01000011_1100_011: DATA = 1'b1;
            15'b01000011_1100_100: DATA = 1'b1;
            15'b01000011_1100_101: DATA = 1'b0;
            15'b01000011_1100_110: DATA = 1'b0;
            15'b01000011_1100_111: DATA = 1'b0;
            // C Row 13
            15'b01000011_1101_000: DATA = 1'b0;
            15'b01000011_1101_001: DATA = 1'b0;
            15'b01000011_1101_010: DATA = 1'b0;
            15'b01000011_1101_011: DATA = 1'b0;
            15'b01000011_1101_100: DATA = 1'b0;
            15'b01000011_1101_101: DATA = 1'b0;
            15'b01000011_1101_110: DATA = 1'b0;
            15'b01000011_1101_111: DATA = 1'b0;
            // C Row 14
            15'b01000011_1110_000: DATA = 1'b0;
            15'b01000011_1110_001: DATA = 1'b0;
            15'b01000011_1110_010: DATA = 1'b0;
            15'b01000011_1110_011: DATA = 1'b0;
            15'b01000011_1110_100: DATA = 1'b0;
            15'b01000011_1110_101: DATA = 1'b0;
            15'b01000011_1110_110: DATA = 1'b0;
            15'b01000011_1110_111: DATA = 1'b0;
            // C Row 15
            15'b01000011_1111_000: DATA = 1'b0;
            15'b01000011_1111_001: DATA = 1'b0;
            15'b01000011_1111_010: DATA = 1'b0;
            15'b01000011_1111_011: DATA = 1'b0;
            15'b01000011_1111_100: DATA = 1'b0;
            15'b01000011_1111_101: DATA = 1'b0;
            15'b01000011_1111_110: DATA = 1'b0;
            15'b01000011_1111_111: DATA = 1'b0;
            // D Row 0
            15'b01000100_0000_000: DATA = 1'b0;
            15'b01000100_0000_001: DATA = 1'b0;
            15'b01000100_0000_010: DATA = 1'b0;
            15'b01000100_0000_011: DATA = 1'b0;
            15'b01000100_0000_100: DATA = 1'b0;
            15'b01000100_0000_101: DATA = 1'b0;
            15'b01000100_0000_110: DATA = 1'b0;
            15'b01000100_0000_111: DATA = 1'b0;
            // D Row 1
            15'b01000100_0001_000: DATA = 1'b0;
            15'b01000100_0001_001: DATA = 1'b0;
            15'b01000100_0001_010: DATA = 1'b0;
            15'b01000100_0001_011: DATA = 1'b0;
            15'b01000100_0001_100: DATA = 1'b0;
            15'b01000100_0001_101: DATA = 1'b0;
            15'b01000100_0001_110: DATA = 1'b0;
            15'b01000100_0001_111: DATA = 1'b0;
            // D Row 2
            15'b01000100_0010_000: DATA = 1'b0;
            15'b01000100_0010_001: DATA = 1'b0;
            15'b01000100_0010_010: DATA = 1'b0;
            15'b01000100_0010_011: DATA = 1'b0;
            15'b01000100_0010_100: DATA = 1'b0;
            15'b01000100_0010_101: DATA = 1'b0;
            15'b01000100_0010_110: DATA = 1'b0;
            15'b01000100_0010_111: DATA = 1'b0;
            // D Row 3
            15'b01000100_0011_000: DATA = 1'b1;
            15'b01000100_0011_001: DATA = 1'b1;
            15'b01000100_0011_010: DATA = 1'b1;
            15'b01000100_0011_011: DATA = 1'b1;
            15'b01000100_0011_100: DATA = 1'b1;
            15'b01000100_0011_101: DATA = 1'b0;
            15'b01000100_0011_110: DATA = 1'b0;
            15'b01000100_0011_111: DATA = 1'b0;
            // D Row 4
            15'b01000100_0100_000: DATA = 1'b1;
            15'b01000100_0100_001: DATA = 1'b1;
            15'b01000100_0100_010: DATA = 1'b0;
            15'b01000100_0100_011: DATA = 1'b0;
            15'b01000100_0100_100: DATA = 1'b1;
            15'b01000100_0100_101: DATA = 1'b1;
            15'b01000100_0100_110: DATA = 1'b0;
            15'b01000100_0100_111: DATA = 1'b0;
            // D Row 5
            15'b01000100_0101_000: DATA = 1'b1;
            15'b01000100_0101_001: DATA = 1'b1;
            15'b01000100_0101_010: DATA = 1'b0;
            15'b01000100_0101_011: DATA = 1'b0;
            15'b01000100_0101_100: DATA = 1'b0;
            15'b01000100_0101_101: DATA = 1'b1;
            15'b01000100_0101_110: DATA = 1'b0;
            15'b01000100_0101_111: DATA = 1'b0;
            // D Row 6
            15'b01000100_0110_000: DATA = 1'b1;
            15'b01000100_0110_001: DATA = 1'b1;
            15'b01000100_0110_010: DATA = 1'b0;
            15'b01000100_0110_011: DATA = 1'b0;
            15'b01000100_0110_100: DATA = 1'b0;
            15'b01000100_0110_101: DATA = 1'b1;
            15'b01000100_0110_110: DATA = 1'b1;
            15'b01000100_0110_111: DATA = 1'b0;
            // D Row 7
            15'b01000100_0111_000: DATA = 1'b1;
            15'b01000100_0111_001: DATA = 1'b1;
            15'b01000100_0111_010: DATA = 1'b0;
            15'b01000100_0111_011: DATA = 1'b0;
            15'b01000100_0111_100: DATA = 1'b0;
            15'b01000100_0111_101: DATA = 1'b1;
            15'b01000100_0111_110: DATA = 1'b1;
            15'b01000100_0111_111: DATA = 1'b0;
            // D Row 8
            15'b01000100_1000_000: DATA = 1'b1;
            15'b01000100_1000_001: DATA = 1'b1;
            15'b01000100_1000_010: DATA = 1'b0;
            15'b01000100_1000_011: DATA = 1'b0;
            15'b01000100_1000_100: DATA = 1'b0;
            15'b01000100_1000_101: DATA = 1'b1;
            15'b01000100_1000_110: DATA = 1'b1;
            15'b01000100_1000_111: DATA = 1'b0;
            // D Row 9
            15'b01000100_1001_000: DATA = 1'b1;
            15'b01000100_1001_001: DATA = 1'b1;
            15'b01000100_1001_010: DATA = 1'b0;
            15'b01000100_1001_011: DATA = 1'b0;
            15'b01000100_1001_100: DATA = 1'b0;
            15'b01000100_1001_101: DATA = 1'b1;
            15'b01000100_1001_110: DATA = 1'b1;
            15'b01000100_1001_111: DATA = 1'b0;
            // D Row 10
            15'b01000100_1010_000: DATA = 1'b1;
            15'b01000100_1010_001: DATA = 1'b1;
            15'b01000100_1010_010: DATA = 1'b0;
            15'b01000100_1010_011: DATA = 1'b0;
            15'b01000100_1010_100: DATA = 1'b1;
            15'b01000100_1010_101: DATA = 1'b0;
            15'b01000100_1010_110: DATA = 1'b0;
            15'b01000100_1010_111: DATA = 1'b0;
            // D Row 11
            15'b01000100_1011_000: DATA = 1'b1;
            15'b01000100_1011_001: DATA = 1'b1;
            15'b01000100_1011_010: DATA = 1'b0;
            15'b01000100_1011_011: DATA = 1'b0;
            15'b01000100_1011_100: DATA = 1'b1;
            15'b01000100_1011_101: DATA = 1'b1;
            15'b01000100_1011_110: DATA = 1'b0;
            15'b01000100_1011_111: DATA = 1'b0;
            // D Row 12
            15'b01000100_1100_000: DATA = 1'b1;
            15'b01000100_1100_001: DATA = 1'b1;
            15'b01000100_1100_010: DATA = 1'b1;
            15'b01000100_1100_011: DATA = 1'b1;
            15'b01000100_1100_100: DATA = 1'b1;
            15'b01000100_1100_101: DATA = 1'b0;
            15'b01000100_1100_110: DATA = 1'b0;
            15'b01000100_1100_111: DATA = 1'b0;
            // D Row 13
            15'b01000100_1101_000: DATA = 1'b0;
            15'b01000100_1101_001: DATA = 1'b0;
            15'b01000100_1101_010: DATA = 1'b0;
            15'b01000100_1101_011: DATA = 1'b0;
            15'b01000100_1101_100: DATA = 1'b0;
            15'b01000100_1101_101: DATA = 1'b0;
            15'b01000100_1101_110: DATA = 1'b0;
            15'b01000100_1101_111: DATA = 1'b0;
            // D Row 14
            15'b01000100_1110_000: DATA = 1'b0;
            15'b01000100_1110_001: DATA = 1'b0;
            15'b01000100_1110_010: DATA = 1'b0;
            15'b01000100_1110_011: DATA = 1'b0;
            15'b01000100_1110_100: DATA = 1'b0;
            15'b01000100_1110_101: DATA = 1'b0;
            15'b01000100_1110_110: DATA = 1'b0;
            15'b01000100_1110_111: DATA = 1'b0;
            // D Row 15
            15'b01000100_1111_000: DATA = 1'b0;
            15'b01000100_1111_001: DATA = 1'b0;
            15'b01000100_1111_010: DATA = 1'b0;
            15'b01000100_1111_011: DATA = 1'b0;
            15'b01000100_1111_100: DATA = 1'b0;
            15'b01000100_1111_101: DATA = 1'b0;
            15'b01000100_1111_110: DATA = 1'b0;
            15'b01000100_1111_111: DATA = 1'b0;
            // E Row 0
            15'b01000101_0000_000: DATA = 1'b0;
            15'b01000101_0000_001: DATA = 1'b0;
            15'b01000101_0000_010: DATA = 1'b0;
            15'b01000101_0000_011: DATA = 1'b0;
            15'b01000101_0000_100: DATA = 1'b0;
            15'b01000101_0000_101: DATA = 1'b0;
            15'b01000101_0000_110: DATA = 1'b0;
            15'b01000101_0000_111: DATA = 1'b0;
            // E Row 1
            15'b01000101_0001_000: DATA = 1'b0;
            15'b01000101_0001_001: DATA = 1'b0;
            15'b01000101_0001_010: DATA = 1'b0;
            15'b01000101_0001_011: DATA = 1'b0;
            15'b01000101_0001_100: DATA = 1'b0;
            15'b01000101_0001_101: DATA = 1'b0;
            15'b01000101_0001_110: DATA = 1'b0;
            15'b01000101_0001_111: DATA = 1'b0;
            // E Row 2
            15'b01000101_0010_000: DATA = 1'b0;
            15'b01000101_0010_001: DATA = 1'b0;
            15'b01000101_0010_010: DATA = 1'b0;
            15'b01000101_0010_011: DATA = 1'b0;
            15'b01000101_0010_100: DATA = 1'b0;
            15'b01000101_0010_101: DATA = 1'b0;
            15'b01000101_0010_110: DATA = 1'b0;
            15'b01000101_0010_111: DATA = 1'b0;
            // E Row 3
            15'b01000101_0011_000: DATA = 1'b1;
            15'b01000101_0011_001: DATA = 1'b1;
            15'b01000101_0011_010: DATA = 1'b1;
            15'b01000101_0011_011: DATA = 1'b1;
            15'b01000101_0011_100: DATA = 1'b1;
            15'b01000101_0011_101: DATA = 1'b1;
            15'b01000101_0011_110: DATA = 1'b1;
            15'b01000101_0011_111: DATA = 1'b0;
            // E Row 4
            15'b01000101_0100_000: DATA = 1'b1;
            15'b01000101_0100_001: DATA = 1'b1;
            15'b01000101_0100_010: DATA = 1'b1;
            15'b01000101_0100_011: DATA = 1'b1;
            15'b01000101_0100_100: DATA = 1'b1;
            15'b01000101_0100_101: DATA = 1'b1;
            15'b01000101_0100_110: DATA = 1'b1;
            15'b01000101_0100_111: DATA = 1'b0;
            // E Row 5
            15'b01000101_0101_000: DATA = 1'b1;
            15'b01000101_0101_001: DATA = 1'b1;
            15'b01000101_0101_010: DATA = 1'b0;
            15'b01000101_0101_011: DATA = 1'b0;
            15'b01000101_0101_100: DATA = 1'b0;
            15'b01000101_0101_101: DATA = 1'b0;
            15'b01000101_0101_110: DATA = 1'b0;
            15'b01000101_0101_111: DATA = 1'b0;
            // E Row 6
            15'b01000101_0110_000: DATA = 1'b1;
            15'b01000101_0110_001: DATA = 1'b1;
            15'b01000101_0110_010: DATA = 1'b0;
            15'b01000101_0110_011: DATA = 1'b0;
            15'b01000101_0110_100: DATA = 1'b0;
            15'b01000101_0110_101: DATA = 1'b0;
            15'b01000101_0110_110: DATA = 1'b0;
            15'b01000101_0110_111: DATA = 1'b0;
            // E Row 7
            15'b01000101_0111_000: DATA = 1'b1;
            15'b01000101_0111_001: DATA = 1'b1;
            15'b01000101_0111_010: DATA = 1'b1;
            15'b01000101_0111_011: DATA = 1'b1;
            15'b01000101_0111_100: DATA = 1'b1;
            15'b01000101_0111_101: DATA = 1'b1;
            15'b01000101_0111_110: DATA = 1'b0;
            15'b01000101_0111_111: DATA = 1'b0;
            // E Row 8
            15'b01000101_1000_000: DATA = 1'b1;
            15'b01000101_1000_001: DATA = 1'b1;
            15'b01000101_1000_010: DATA = 1'b1;
            15'b01000101_1000_011: DATA = 1'b1;
            15'b01000101_1000_100: DATA = 1'b1;
            15'b01000101_1000_101: DATA = 1'b1;
            15'b01000101_1000_110: DATA = 1'b0;
            15'b01000101_1000_111: DATA = 1'b0;
            // E Row 9
            15'b01000101_1001_000: DATA = 1'b1;
            15'b01000101_1001_001: DATA = 1'b1;
            15'b01000101_1001_010: DATA = 1'b0;
            15'b01000101_1001_011: DATA = 1'b0;
            15'b01000101_1001_100: DATA = 1'b0;
            15'b01000101_1001_101: DATA = 1'b0;
            15'b01000101_1001_110: DATA = 1'b0;
            15'b01000101_1001_111: DATA = 1'b0;
            // E Row 10
            15'b01000101_1010_000: DATA = 1'b1;
            15'b01000101_1010_001: DATA = 1'b1;
            15'b01000101_1010_010: DATA = 1'b0;
            15'b01000101_1010_011: DATA = 1'b0;
            15'b01000101_1010_100: DATA = 1'b0;
            15'b01000101_1010_101: DATA = 1'b0;
            15'b01000101_1010_110: DATA = 1'b0;
            15'b01000101_1010_111: DATA = 1'b0;
            // E Row 11
            15'b01000101_1011_000: DATA = 1'b1;
            15'b01000101_1011_001: DATA = 1'b1;
            15'b01000101_1011_010: DATA = 1'b1;
            15'b01000101_1011_011: DATA = 1'b1;
            15'b01000101_1011_100: DATA = 1'b1;
            15'b01000101_1011_101: DATA = 1'b1;
            15'b01000101_1011_110: DATA = 1'b1;
            15'b01000101_1011_111: DATA = 1'b0;
            // E Row 12
            15'b01000101_1100_000: DATA = 1'b1;
            15'b01000101_1100_001: DATA = 1'b1;
            15'b01000101_1100_010: DATA = 1'b1;
            15'b01000101_1100_011: DATA = 1'b1;
            15'b01000101_1100_100: DATA = 1'b1;
            15'b01000101_1100_101: DATA = 1'b1;
            15'b01000101_1100_110: DATA = 1'b1;
            15'b01000101_1100_111: DATA = 1'b0;
            // E Row 13
            15'b01000101_1101_000: DATA = 1'b0;
            15'b01000101_1101_001: DATA = 1'b0;
            15'b01000101_1101_010: DATA = 1'b0;
            15'b01000101_1101_011: DATA = 1'b0;
            15'b01000101_1101_100: DATA = 1'b0;
            15'b01000101_1101_101: DATA = 1'b0;
            15'b01000101_1101_110: DATA = 1'b0;
            15'b01000101_1101_111: DATA = 1'b0;
            // E Row 14
            15'b01000101_1110_000: DATA = 1'b0;
            15'b01000101_1110_001: DATA = 1'b0;
            15'b01000101_1110_010: DATA = 1'b0;
            15'b01000101_1110_011: DATA = 1'b0;
            15'b01000101_1110_100: DATA = 1'b0;
            15'b01000101_1110_101: DATA = 1'b0;
            15'b01000101_1110_110: DATA = 1'b0;
            15'b01000101_1110_111: DATA = 1'b0;
            // E Row 15
            15'b01000101_1111_000: DATA = 1'b0;
            15'b01000101_1111_001: DATA = 1'b0;
            15'b01000101_1111_010: DATA = 1'b0;
            15'b01000101_1111_011: DATA = 1'b0;
            15'b01000101_1111_100: DATA = 1'b0;
            15'b01000101_1111_101: DATA = 1'b0;
            15'b01000101_1111_110: DATA = 1'b0;
            15'b01000101_1111_111: DATA = 1'b0;
            // F Row 0
            15'b01000110_0000_000: DATA = 1'b0;
            15'b01000110_0000_001: DATA = 1'b0;
            15'b01000110_0000_010: DATA = 1'b0;
            15'b01000110_0000_011: DATA = 1'b0;
            15'b01000110_0000_100: DATA = 1'b0;
            15'b01000110_0000_101: DATA = 1'b0;
            15'b01000110_0000_110: DATA = 1'b0;
            15'b01000110_0000_111: DATA = 1'b0;
            // F Row 1
            15'b01000110_0001_000: DATA = 1'b0;
            15'b01000110_0001_001: DATA = 1'b0;
            15'b01000110_0001_010: DATA = 1'b0;
            15'b01000110_0001_011: DATA = 1'b0;
            15'b01000110_0001_100: DATA = 1'b0;
            15'b01000110_0001_101: DATA = 1'b0;
            15'b01000110_0001_110: DATA = 1'b0;
            15'b01000110_0001_111: DATA = 1'b0;
            // F Row 2
            15'b01000110_0010_000: DATA = 1'b0;
            15'b01000110_0010_001: DATA = 1'b0;
            15'b01000110_0010_010: DATA = 1'b0;
            15'b01000110_0010_011: DATA = 1'b0;
            15'b01000110_0010_100: DATA = 1'b0;
            15'b01000110_0010_101: DATA = 1'b0;
            15'b01000110_0010_110: DATA = 1'b0;
            15'b01000110_0010_111: DATA = 1'b0;
            // F Row 3
            15'b01000110_0011_000: DATA = 1'b1;
            15'b01000110_0011_001: DATA = 1'b1;
            15'b01000110_0011_010: DATA = 1'b1;
            15'b01000110_0011_011: DATA = 1'b1;
            15'b01000110_0011_100: DATA = 1'b1;
            15'b01000110_0011_101: DATA = 1'b1;
            15'b01000110_0011_110: DATA = 1'b1;
            15'b01000110_0011_111: DATA = 1'b0;
            // F Row 4
            15'b01000110_0100_000: DATA = 1'b1;
            15'b01000110_0100_001: DATA = 1'b1;
            15'b01000110_0100_010: DATA = 1'b1;
            15'b01000110_0100_011: DATA = 1'b1;
            15'b01000110_0100_100: DATA = 1'b1;
            15'b01000110_0100_101: DATA = 1'b1;
            15'b01000110_0100_110: DATA = 1'b1;
            15'b01000110_0100_111: DATA = 1'b0;
            // F Row 5
            15'b01000110_0101_000: DATA = 1'b1;
            15'b01000110_0101_001: DATA = 1'b1;
            15'b01000110_0101_010: DATA = 1'b0;
            15'b01000110_0101_011: DATA = 1'b0;
            15'b01000110_0101_100: DATA = 1'b0;
            15'b01000110_0101_101: DATA = 1'b0;
            15'b01000110_0101_110: DATA = 1'b0;
            15'b01000110_0101_111: DATA = 1'b0;
            // F Row 6
            15'b01000110_0110_000: DATA = 1'b1;
            15'b01000110_0110_001: DATA = 1'b1;
            15'b01000110_0110_010: DATA = 1'b0;
            15'b01000110_0110_011: DATA = 1'b0;
            15'b01000110_0110_100: DATA = 1'b0;
            15'b01000110_0110_101: DATA = 1'b0;
            15'b01000110_0110_110: DATA = 1'b0;
            15'b01000110_0110_111: DATA = 1'b0;
            // F Row 7
            15'b01000110_0111_000: DATA = 1'b1;
            15'b01000110_0111_001: DATA = 1'b1;
            15'b01000110_0111_010: DATA = 1'b1;
            15'b01000110_0111_011: DATA = 1'b1;
            15'b01000110_0111_100: DATA = 1'b1;
            15'b01000110_0111_101: DATA = 1'b1;
            15'b01000110_0111_110: DATA = 1'b0;
            15'b01000110_0111_111: DATA = 1'b0;
            // F Row 8
            15'b01000110_1000_000: DATA = 1'b1;
            15'b01000110_1000_001: DATA = 1'b1;
            15'b01000110_1000_010: DATA = 1'b1;
            15'b01000110_1000_011: DATA = 1'b1;
            15'b01000110_1000_100: DATA = 1'b1;
            15'b01000110_1000_101: DATA = 1'b1;
            15'b01000110_1000_110: DATA = 1'b0;
            15'b01000110_1000_111: DATA = 1'b0;
            // F Row 9
            15'b01000110_1001_000: DATA = 1'b1;
            15'b01000110_1001_001: DATA = 1'b1;
            15'b01000110_1001_010: DATA = 1'b0;
            15'b01000110_1001_011: DATA = 1'b0;
            15'b01000110_1001_100: DATA = 1'b0;
            15'b01000110_1001_101: DATA = 1'b0;
            15'b01000110_1001_110: DATA = 1'b0;
            15'b01000110_1001_111: DATA = 1'b0;
            // F Row 10
            15'b01000110_1010_000: DATA = 1'b1;
            15'b01000110_1010_001: DATA = 1'b1;
            15'b01000110_1010_010: DATA = 1'b0;
            15'b01000110_1010_011: DATA = 1'b0;
            15'b01000110_1010_100: DATA = 1'b0;
            15'b01000110_1010_101: DATA = 1'b0;
            15'b01000110_1010_110: DATA = 1'b0;
            15'b01000110_1010_111: DATA = 1'b0;
            // F Row 11
            15'b01000110_1011_000: DATA = 1'b1;
            15'b01000110_1011_001: DATA = 1'b1;
            15'b01000110_1011_010: DATA = 1'b0;
            15'b01000110_1011_011: DATA = 1'b0;
            15'b01000110_1011_100: DATA = 1'b0;
            15'b01000110_1011_101: DATA = 1'b0;
            15'b01000110_1011_110: DATA = 1'b0;
            15'b01000110_1011_111: DATA = 1'b0;
            // F Row 12
            15'b01000110_1100_000: DATA = 1'b1;
            15'b01000110_1100_001: DATA = 1'b1;
            15'b01000110_1100_010: DATA = 1'b0;
            15'b01000110_1100_011: DATA = 1'b0;
            15'b01000110_1100_100: DATA = 1'b0;
            15'b01000110_1100_101: DATA = 1'b0;
            15'b01000110_1100_110: DATA = 1'b0;
            15'b01000110_1100_111: DATA = 1'b0;
            // F Row 13
            15'b01000110_1101_000: DATA = 1'b0;
            15'b01000110_1101_001: DATA = 1'b0;
            15'b01000110_1101_010: DATA = 1'b0;
            15'b01000110_1101_011: DATA = 1'b0;
            15'b01000110_1101_100: DATA = 1'b0;
            15'b01000110_1101_101: DATA = 1'b0;
            15'b01000110_1101_110: DATA = 1'b0;
            15'b01000110_1101_111: DATA = 1'b0;
            // F Row 14
            15'b01000110_1110_000: DATA = 1'b0;
            15'b01000110_1110_001: DATA = 1'b0;
            15'b01000110_1110_010: DATA = 1'b0;
            15'b01000110_1110_011: DATA = 1'b0;
            15'b01000110_1110_100: DATA = 1'b0;
            15'b01000110_1110_101: DATA = 1'b0;
            15'b01000110_1110_110: DATA = 1'b0;
            15'b01000110_1110_111: DATA = 1'b0;
            // F Row 15
            15'b01000110_1111_000: DATA = 1'b0;
            15'b01000110_1111_001: DATA = 1'b0;
            15'b01000110_1111_010: DATA = 1'b0;
            15'b01000110_1111_011: DATA = 1'b0;
            15'b01000110_1111_100: DATA = 1'b0;
            15'b01000110_1111_101: DATA = 1'b0;
            15'b01000110_1111_110: DATA = 1'b0;
            15'b01000110_1111_111: DATA = 1'b0;
            // G Row 0
            15'b01000111_0000_000: DATA = 1'b0;
            15'b01000111_0000_001: DATA = 1'b0;
            15'b01000111_0000_010: DATA = 1'b0;
            15'b01000111_0000_011: DATA = 1'b0;
            15'b01000111_0000_100: DATA = 1'b0;
            15'b01000111_0000_101: DATA = 1'b0;
            15'b01000111_0000_110: DATA = 1'b0;
            15'b01000111_0000_111: DATA = 1'b0;
            // G Row 1
            15'b01000111_0001_000: DATA = 1'b0;
            15'b01000111_0001_001: DATA = 1'b0;
            15'b01000111_0001_010: DATA = 1'b0;
            15'b01000111_0001_011: DATA = 1'b0;
            15'b01000111_0001_100: DATA = 1'b0;
            15'b01000111_0001_101: DATA = 1'b0;
            15'b01000111_0001_110: DATA = 1'b0;
            15'b01000111_0001_111: DATA = 1'b0;
            // G Row 2
            15'b01000111_0010_000: DATA = 1'b0;
            15'b01000111_0010_001: DATA = 1'b0;
            15'b01000111_0010_010: DATA = 1'b0;
            15'b01000111_0010_011: DATA = 1'b0;
            15'b01000111_0010_100: DATA = 1'b0;
            15'b01000111_0010_101: DATA = 1'b0;
            15'b01000111_0010_110: DATA = 1'b0;
            15'b01000111_0010_111: DATA = 1'b0;
            // G Row 3
            15'b01000111_0011_000: DATA = 1'b0;
            15'b01000111_0011_001: DATA = 1'b0;
            15'b01000111_0011_010: DATA = 1'b1;
            15'b01000111_0011_011: DATA = 1'b1;
            15'b01000111_0011_100: DATA = 1'b1;
            15'b01000111_0011_101: DATA = 1'b0;
            15'b01000111_0011_110: DATA = 1'b0;
            15'b01000111_0011_111: DATA = 1'b0;
            // G Row 4
            15'b01000111_0100_000: DATA = 1'b0;
            15'b01000111_0100_001: DATA = 1'b1;
            15'b01000111_0100_010: DATA = 1'b1;
            15'b01000111_0100_011: DATA = 1'b1;
            15'b01000111_0100_100: DATA = 1'b1;
            15'b01000111_0100_101: DATA = 1'b1;
            15'b01000111_0100_110: DATA = 1'b0;
            15'b01000111_0100_111: DATA = 1'b0;
            // G Row 5
            15'b01000111_0101_000: DATA = 1'b1;
            15'b01000111_0101_001: DATA = 1'b1;
            15'b01000111_0101_010: DATA = 1'b0;
            15'b01000111_0101_011: DATA = 1'b0;
            15'b01000111_0101_100: DATA = 1'b0;
            15'b01000111_0101_101: DATA = 1'b1;
            15'b01000111_0101_110: DATA = 1'b1;
            15'b01000111_0101_111: DATA = 1'b0;
            // G Row 6
            15'b01000111_0110_000: DATA = 1'b1;
            15'b01000111_0110_001: DATA = 1'b1;
            15'b01000111_0110_010: DATA = 1'b0;
            15'b01000111_0110_011: DATA = 1'b0;
            15'b01000111_0110_100: DATA = 1'b0;
            15'b01000111_0110_101: DATA = 1'b0;
            15'b01000111_0110_110: DATA = 1'b0;
            15'b01000111_0110_111: DATA = 1'b0;
            // G Row 7
            15'b01000111_0111_000: DATA = 1'b1;
            15'b01000111_0111_001: DATA = 1'b1;
            15'b01000111_0111_010: DATA = 1'b0;
            15'b01000111_0111_011: DATA = 1'b0;
            15'b01000111_0111_100: DATA = 1'b0;
            15'b01000111_0111_101: DATA = 1'b0;
            15'b01000111_0111_110: DATA = 1'b0;
            15'b01000111_0111_111: DATA = 1'b0;
            // G Row 8
            15'b01000111_1000_000: DATA = 1'b1;
            15'b01000111_1000_001: DATA = 1'b1;
            15'b01000111_1000_010: DATA = 1'b0;
            15'b01000111_1000_011: DATA = 1'b1;
            15'b01000111_1000_100: DATA = 1'b1;
            15'b01000111_1000_101: DATA = 1'b1;
            15'b01000111_1000_110: DATA = 1'b1;
            15'b01000111_1000_111: DATA = 1'b0;
            // G Row 9
            15'b01000111_1001_000: DATA = 1'b1;
            15'b01000111_1001_001: DATA = 1'b1;
            15'b01000111_1001_010: DATA = 1'b0;
            15'b01000111_1001_011: DATA = 1'b0;
            15'b01000111_1001_100: DATA = 1'b0;
            15'b01000111_1001_101: DATA = 1'b1;
            15'b01000111_1001_110: DATA = 1'b1;
            15'b01000111_1001_111: DATA = 1'b0;
            // G Row 10
            15'b01000111_1010_000: DATA = 1'b1;
            15'b01000111_1010_001: DATA = 1'b1;
            15'b01000111_1010_010: DATA = 1'b0;
            15'b01000111_1010_011: DATA = 1'b0;
            15'b01000111_1010_100: DATA = 1'b0;
            15'b01000111_1010_101: DATA = 1'b1;
            15'b01000111_1010_110: DATA = 1'b1;
            15'b01000111_1010_111: DATA = 1'b0;
            // G Row 11
            15'b01000111_1011_000: DATA = 1'b0;
            15'b01000111_1011_001: DATA = 1'b1;
            15'b01000111_1011_010: DATA = 1'b1;
            15'b01000111_1011_011: DATA = 1'b1;
            15'b01000111_1011_100: DATA = 1'b1;
            15'b01000111_1011_101: DATA = 1'b1;
            15'b01000111_1011_110: DATA = 1'b0;
            15'b01000111_1011_111: DATA = 1'b0;
            // G Row 12
            15'b01000111_1100_000: DATA = 1'b0;
            15'b01000111_1100_001: DATA = 1'b0;
            15'b01000111_1100_010: DATA = 1'b1;
            15'b01000111_1100_011: DATA = 1'b1;
            15'b01000111_1100_100: DATA = 1'b1;
            15'b01000111_1100_101: DATA = 1'b0;
            15'b01000111_1100_110: DATA = 1'b0;
            15'b01000111_1100_111: DATA = 1'b0;
            // G Row 13
            15'b01000111_1101_000: DATA = 1'b0;
            15'b01000111_1101_001: DATA = 1'b0;
            15'b01000111_1101_010: DATA = 1'b0;
            15'b01000111_1101_011: DATA = 1'b0;
            15'b01000111_1101_100: DATA = 1'b0;
            15'b01000111_1101_101: DATA = 1'b0;
            15'b01000111_1101_110: DATA = 1'b0;
            15'b01000111_1101_111: DATA = 1'b0;
            // G Row 14
            15'b01000111_1110_000: DATA = 1'b0;
            15'b01000111_1110_001: DATA = 1'b0;
            15'b01000111_1110_010: DATA = 1'b0;
            15'b01000111_1110_011: DATA = 1'b0;
            15'b01000111_1110_100: DATA = 1'b0;
            15'b01000111_1110_101: DATA = 1'b0;
            15'b01000111_1110_110: DATA = 1'b0;
            15'b01000111_1110_111: DATA = 1'b0;
            // G Row 15
            15'b01000111_1111_000: DATA = 1'b0;
            15'b01000111_1111_001: DATA = 1'b0;
            15'b01000111_1111_010: DATA = 1'b0;
            15'b01000111_1111_011: DATA = 1'b0;
            15'b01000111_1111_100: DATA = 1'b0;
            15'b01000111_1111_101: DATA = 1'b0;
            15'b01000111_1111_110: DATA = 1'b0;
            15'b01000111_1111_111: DATA = 1'b0;
            // H Row 0
            15'b01001000_0000_000: DATA = 1'b0;
            15'b01001000_0000_001: DATA = 1'b0;
            15'b01001000_0000_010: DATA = 1'b0;
            15'b01001000_0000_011: DATA = 1'b0;
            15'b01001000_0000_100: DATA = 1'b0;
            15'b01001000_0000_101: DATA = 1'b0;
            15'b01001000_0000_110: DATA = 1'b0;
            15'b01001000_0000_111: DATA = 1'b0;
            // H Row 1
            15'b01001000_0001_000: DATA = 1'b0;
            15'b01001000_0001_001: DATA = 1'b0;
            15'b01001000_0001_010: DATA = 1'b0;
            15'b01001000_0001_011: DATA = 1'b0;
            15'b01001000_0001_100: DATA = 1'b0;
            15'b01001000_0001_101: DATA = 1'b0;
            15'b01001000_0001_110: DATA = 1'b0;
            15'b01001000_0001_111: DATA = 1'b0;
            // H Row 2
            15'b01001000_0010_000: DATA = 1'b0;
            15'b01001000_0010_001: DATA = 1'b0;
            15'b01001000_0010_010: DATA = 1'b0;
            15'b01001000_0010_011: DATA = 1'b0;
            15'b01001000_0010_100: DATA = 1'b0;
            15'b01001000_0010_101: DATA = 1'b0;
            15'b01001000_0010_110: DATA = 1'b0;
            15'b01001000_0010_111: DATA = 1'b0;
            // H Row 3
            15'b01001000_0011_000: DATA = 1'b1;
            15'b01001000_0011_001: DATA = 1'b1;
            15'b01001000_0011_010: DATA = 1'b0;
            15'b01001000_0011_011: DATA = 1'b0;
            15'b01001000_0011_100: DATA = 1'b0;
            15'b01001000_0011_101: DATA = 1'b1;
            15'b01001000_0011_110: DATA = 1'b1;
            15'b01001000_0011_111: DATA = 1'b0;
            // H Row 4
            15'b01001000_0100_000: DATA = 1'b1;
            15'b01001000_0100_001: DATA = 1'b1;
            15'b01001000_0100_010: DATA = 1'b0;
            15'b01001000_0100_011: DATA = 1'b0;
            15'b01001000_0100_100: DATA = 1'b0;
            15'b01001000_0100_101: DATA = 1'b1;
            15'b01001000_0100_110: DATA = 1'b1;
            15'b01001000_0100_111: DATA = 1'b0;
            // H Row 5
            15'b01001000_0101_000: DATA = 1'b1;
            15'b01001000_0101_001: DATA = 1'b1;
            15'b01001000_0101_010: DATA = 1'b0;
            15'b01001000_0101_011: DATA = 1'b0;
            15'b01001000_0101_100: DATA = 1'b0;
            15'b01001000_0101_101: DATA = 1'b1;
            15'b01001000_0101_110: DATA = 1'b1;
            15'b01001000_0101_111: DATA = 1'b0;
            // H Row 6
            15'b01001000_0110_000: DATA = 1'b1;
            15'b01001000_0110_001: DATA = 1'b1;
            15'b01001000_0110_010: DATA = 1'b0;
            15'b01001000_0110_011: DATA = 1'b0;
            15'b01001000_0110_100: DATA = 1'b0;
            15'b01001000_0110_101: DATA = 1'b1;
            15'b01001000_0110_110: DATA = 1'b1;
            15'b01001000_0110_111: DATA = 1'b0;
            // H Row 7
            15'b01001000_0111_000: DATA = 1'b1;
            15'b01001000_0111_001: DATA = 1'b1;
            15'b01001000_0111_010: DATA = 1'b1;
            15'b01001000_0111_011: DATA = 1'b1;
            15'b01001000_0111_100: DATA = 1'b1;
            15'b01001000_0111_101: DATA = 1'b1;
            15'b01001000_0111_110: DATA = 1'b1;
            15'b01001000_0111_111: DATA = 1'b0;
            // H Row 8
            15'b01001000_1000_000: DATA = 1'b1;
            15'b01001000_1000_001: DATA = 1'b1;
            15'b01001000_1000_010: DATA = 1'b1;
            15'b01001000_1000_011: DATA = 1'b1;
            15'b01001000_1000_100: DATA = 1'b1;
            15'b01001000_1000_101: DATA = 1'b1;
            15'b01001000_1000_110: DATA = 1'b1;
            15'b01001000_1000_111: DATA = 1'b0;
            // H Row 9
            15'b01001000_1001_000: DATA = 1'b1;
            15'b01001000_1001_001: DATA = 1'b1;
            15'b01001000_1001_010: DATA = 1'b0;
            15'b01001000_1001_011: DATA = 1'b0;
            15'b01001000_1001_100: DATA = 1'b0;
            15'b01001000_1001_101: DATA = 1'b1;
            15'b01001000_1001_110: DATA = 1'b1;
            15'b01001000_1001_111: DATA = 1'b0;
            // H Row 10
            15'b01001000_1010_000: DATA = 1'b1;
            15'b01001000_1010_001: DATA = 1'b1;
            15'b01001000_1010_010: DATA = 1'b0;
            15'b01001000_1010_011: DATA = 1'b0;
            15'b01001000_1010_100: DATA = 1'b0;
            15'b01001000_1010_101: DATA = 1'b1;
            15'b01001000_1010_110: DATA = 1'b1;
            15'b01001000_1010_111: DATA = 1'b0;
            // H Row 11
            15'b01001000_1011_000: DATA = 1'b1;
            15'b01001000_1011_001: DATA = 1'b1;
            15'b01001000_1011_010: DATA = 1'b0;
            15'b01001000_1011_011: DATA = 1'b0;
            15'b01001000_1011_100: DATA = 1'b0;
            15'b01001000_1011_101: DATA = 1'b1;
            15'b01001000_1011_110: DATA = 1'b1;
            15'b01001000_1011_111: DATA = 1'b0;
            // H Row 12
            15'b01001000_1100_000: DATA = 1'b1;
            15'b01001000_1100_001: DATA = 1'b1;
            15'b01001000_1100_010: DATA = 1'b0;
            15'b01001000_1100_011: DATA = 1'b0;
            15'b01001000_1100_100: DATA = 1'b0;
            15'b01001000_1100_101: DATA = 1'b1;
            15'b01001000_1100_110: DATA = 1'b1;
            15'b01001000_1100_111: DATA = 1'b0;
            // H Row 13
            15'b01001000_1101_000: DATA = 1'b0;
            15'b01001000_1101_001: DATA = 1'b0;
            15'b01001000_1101_010: DATA = 1'b0;
            15'b01001000_1101_011: DATA = 1'b0;
            15'b01001000_1101_100: DATA = 1'b0;
            15'b01001000_1101_101: DATA = 1'b0;
            15'b01001000_1101_110: DATA = 1'b0;
            15'b01001000_1101_111: DATA = 1'b0;
            // H Row 14
            15'b01001000_1110_000: DATA = 1'b0;
            15'b01001000_1110_001: DATA = 1'b0;
            15'b01001000_1110_010: DATA = 1'b0;
            15'b01001000_1110_011: DATA = 1'b0;
            15'b01001000_1110_100: DATA = 1'b0;
            15'b01001000_1110_101: DATA = 1'b0;
            15'b01001000_1110_110: DATA = 1'b0;
            15'b01001000_1110_111: DATA = 1'b0;
            // H Row 15
            15'b01001000_1111_000: DATA = 1'b0;
            15'b01001000_1111_001: DATA = 1'b0;
            15'b01001000_1111_010: DATA = 1'b0;
            15'b01001000_1111_011: DATA = 1'b0;
            15'b01001000_1111_100: DATA = 1'b0;
            15'b01001000_1111_101: DATA = 1'b0;
            15'b01001000_1111_110: DATA = 1'b0;
            15'b01001000_1111_111: DATA = 1'b0;
            // I Row 0
            15'b01001001_0000_000: DATA = 1'b0;
            15'b01001001_0000_001: DATA = 1'b0;
            15'b01001001_0000_010: DATA = 1'b0;
            15'b01001001_0000_011: DATA = 1'b0;
            15'b01001001_0000_100: DATA = 1'b0;
            15'b01001001_0000_101: DATA = 1'b0;
            15'b01001001_0000_110: DATA = 1'b0;
            15'b01001001_0000_111: DATA = 1'b0;
            // I Row 1
            15'b01001001_0001_000: DATA = 1'b0;
            15'b01001001_0001_001: DATA = 1'b0;
            15'b01001001_0001_010: DATA = 1'b0;
            15'b01001001_0001_011: DATA = 1'b0;
            15'b01001001_0001_100: DATA = 1'b0;
            15'b01001001_0001_101: DATA = 1'b0;
            15'b01001001_0001_110: DATA = 1'b0;
            15'b01001001_0001_111: DATA = 1'b0;
            // I Row 2
            15'b01001001_0010_000: DATA = 1'b0;
            15'b01001001_0010_001: DATA = 1'b0;
            15'b01001001_0010_010: DATA = 1'b0;
            15'b01001001_0010_011: DATA = 1'b0;
            15'b01001001_0010_100: DATA = 1'b0;
            15'b01001001_0010_101: DATA = 1'b0;
            15'b01001001_0010_110: DATA = 1'b0;
            15'b01001001_0010_111: DATA = 1'b0;
            // I Row 3
            15'b01001001_0011_000: DATA = 1'b1;
            15'b01001001_0011_001: DATA = 1'b1;
            15'b01001001_0011_010: DATA = 1'b1;
            15'b01001001_0011_011: DATA = 1'b1;
            15'b01001001_0011_100: DATA = 1'b1;
            15'b01001001_0011_101: DATA = 1'b1;
            15'b01001001_0011_110: DATA = 1'b1;
            15'b01001001_0011_111: DATA = 1'b0;
            // I Row 4
            15'b01001001_0100_000: DATA = 1'b1;
            15'b01001001_0100_001: DATA = 1'b1;
            15'b01001001_0100_010: DATA = 1'b1;
            15'b01001001_0100_011: DATA = 1'b1;
            15'b01001001_0100_100: DATA = 1'b1;
            15'b01001001_0100_101: DATA = 1'b1;
            15'b01001001_0100_110: DATA = 1'b1;
            15'b01001001_0100_111: DATA = 1'b0;
            // I Row 5
            15'b01001001_0101_000: DATA = 1'b0;
            15'b01001001_0101_001: DATA = 1'b0;
            15'b01001001_0101_010: DATA = 1'b1;
            15'b01001001_0101_011: DATA = 1'b1;
            15'b01001001_0101_100: DATA = 1'b1;
            15'b01001001_0101_101: DATA = 1'b0;
            15'b01001001_0101_110: DATA = 1'b0;
            15'b01001001_0101_111: DATA = 1'b0;
            // I Row 6
            15'b01001001_0110_000: DATA = 1'b0;
            15'b01001001_0110_001: DATA = 1'b0;
            15'b01001001_0110_010: DATA = 1'b1;
            15'b01001001_0110_011: DATA = 1'b1;
            15'b01001001_0110_100: DATA = 1'b1;
            15'b01001001_0110_101: DATA = 1'b0;
            15'b01001001_0110_110: DATA = 1'b0;
            15'b01001001_0110_111: DATA = 1'b0;
            // I Row 7
            15'b01001001_0111_000: DATA = 1'b0;
            15'b01001001_0111_001: DATA = 1'b0;
            15'b01001001_0111_010: DATA = 1'b1;
            15'b01001001_0111_011: DATA = 1'b1;
            15'b01001001_0111_100: DATA = 1'b1;
            15'b01001001_0111_101: DATA = 1'b0;
            15'b01001001_0111_110: DATA = 1'b0;
            15'b01001001_0111_111: DATA = 1'b0;
            // I Row 8
            15'b01001001_1000_000: DATA = 1'b0;
            15'b01001001_1000_001: DATA = 1'b0;
            15'b01001001_1000_010: DATA = 1'b1;
            15'b01001001_1000_011: DATA = 1'b1;
            15'b01001001_1000_100: DATA = 1'b1;
            15'b01001001_1000_101: DATA = 1'b0;
            15'b01001001_1000_110: DATA = 1'b0;
            15'b01001001_1000_111: DATA = 1'b0;
            // I Row 9
            15'b01001001_1001_000: DATA = 1'b0;
            15'b01001001_1001_001: DATA = 1'b0;
            15'b01001001_1001_010: DATA = 1'b1;
            15'b01001001_1001_011: DATA = 1'b1;
            15'b01001001_1001_100: DATA = 1'b1;
            15'b01001001_1001_101: DATA = 1'b0;
            15'b01001001_1001_110: DATA = 1'b0;
            15'b01001001_1001_111: DATA = 1'b0;
            // I Row 10
            15'b01001001_1010_000: DATA = 1'b0;
            15'b01001001_1010_001: DATA = 1'b0;
            15'b01001001_1010_010: DATA = 1'b1;
            15'b01001001_1010_011: DATA = 1'b1;
            15'b01001001_1010_100: DATA = 1'b1;
            15'b01001001_1010_101: DATA = 1'b0;
            15'b01001001_1010_110: DATA = 1'b0;
            15'b01001001_1010_111: DATA = 1'b0;
            // I Row 11
            15'b01001001_1011_000: DATA = 1'b1;
            15'b01001001_1011_001: DATA = 1'b1;
            15'b01001001_1011_010: DATA = 1'b1;
            15'b01001001_1011_011: DATA = 1'b1;
            15'b01001001_1011_100: DATA = 1'b1;
            15'b01001001_1011_101: DATA = 1'b1;
            15'b01001001_1011_110: DATA = 1'b1;
            15'b01001001_1011_111: DATA = 1'b0;
            // I Row 12
            15'b01001001_1100_000: DATA = 1'b1;
            15'b01001001_1100_001: DATA = 1'b1;
            15'b01001001_1100_010: DATA = 1'b1;
            15'b01001001_1100_011: DATA = 1'b1;
            15'b01001001_1100_100: DATA = 1'b1;
            15'b01001001_1100_101: DATA = 1'b1;
            15'b01001001_1100_110: DATA = 1'b1;
            15'b01001001_1100_111: DATA = 1'b0;
            // I Row 13
            15'b01001001_1101_000: DATA = 1'b0;
            15'b01001001_1101_001: DATA = 1'b0;
            15'b01001001_1101_010: DATA = 1'b0;
            15'b01001001_1101_011: DATA = 1'b0;
            15'b01001001_1101_100: DATA = 1'b0;
            15'b01001001_1101_101: DATA = 1'b0;
            15'b01001001_1101_110: DATA = 1'b0;
            15'b01001001_1101_111: DATA = 1'b0;
            // I Row 14
            15'b01001001_1110_000: DATA = 1'b0;
            15'b01001001_1110_001: DATA = 1'b0;
            15'b01001001_1110_010: DATA = 1'b0;
            15'b01001001_1110_011: DATA = 1'b0;
            15'b01001001_1110_100: DATA = 1'b0;
            15'b01001001_1110_101: DATA = 1'b0;
            15'b01001001_1110_110: DATA = 1'b0;
            15'b01001001_1110_111: DATA = 1'b0;
            // I Row 15
            15'b01001001_1111_000: DATA = 1'b0;
            15'b01001001_1111_001: DATA = 1'b0;
            15'b01001001_1111_010: DATA = 1'b0;
            15'b01001001_1111_011: DATA = 1'b0;
            15'b01001001_1111_100: DATA = 1'b0;
            15'b01001001_1111_101: DATA = 1'b0;
            15'b01001001_1111_110: DATA = 1'b0;
            15'b01001001_1111_111: DATA = 1'b0;
            // J Row 0
            15'b01001010_0000_000: DATA = 1'b0;
            15'b01001010_0000_001: DATA = 1'b0;
            15'b01001010_0000_010: DATA = 1'b0;
            15'b01001010_0000_011: DATA = 1'b0;
            15'b01001010_0000_100: DATA = 1'b0;
            15'b01001010_0000_101: DATA = 1'b0;
            15'b01001010_0000_110: DATA = 1'b0;
            15'b01001010_0000_111: DATA = 1'b0;
            // J Row 1
            15'b01001010_0001_000: DATA = 1'b0;
            15'b01001010_0001_001: DATA = 1'b0;
            15'b01001010_0001_010: DATA = 1'b0;
            15'b01001010_0001_011: DATA = 1'b0;
            15'b01001010_0001_100: DATA = 1'b0;
            15'b01001010_0001_101: DATA = 1'b0;
            15'b01001010_0001_110: DATA = 1'b0;
            15'b01001010_0001_111: DATA = 1'b0;
            // J Row 2
            15'b01001010_0010_000: DATA = 1'b0;
            15'b01001010_0010_001: DATA = 1'b0;
            15'b01001010_0010_010: DATA = 1'b0;
            15'b01001010_0010_011: DATA = 1'b0;
            15'b01001010_0010_100: DATA = 1'b0;
            15'b01001010_0010_101: DATA = 1'b0;
            15'b01001010_0010_110: DATA = 1'b0;
            15'b01001010_0010_111: DATA = 1'b0;
            // J Row 3
            15'b01001010_0011_000: DATA = 1'b1;
            15'b01001010_0011_001: DATA = 1'b1;
            15'b01001010_0011_010: DATA = 1'b1;
            15'b01001010_0011_011: DATA = 1'b1;
            15'b01001010_0011_100: DATA = 1'b1;
            15'b01001010_0011_101: DATA = 1'b1;
            15'b01001010_0011_110: DATA = 1'b1;
            15'b01001010_0011_111: DATA = 1'b0;
            // J Row 4
            15'b01001010_0100_000: DATA = 1'b1;
            15'b01001010_0100_001: DATA = 1'b1;
            15'b01001010_0100_010: DATA = 1'b1;
            15'b01001010_0100_011: DATA = 1'b1;
            15'b01001010_0100_100: DATA = 1'b1;
            15'b01001010_0100_101: DATA = 1'b1;
            15'b01001010_0100_110: DATA = 1'b1;
            15'b01001010_0100_111: DATA = 1'b0;
            // J Row 5
            15'b01001010_0101_000: DATA = 1'b0;
            15'b01001010_0101_001: DATA = 1'b0;
            15'b01001010_0101_010: DATA = 1'b0;
            15'b01001010_0101_011: DATA = 1'b0;
            15'b01001010_0101_100: DATA = 1'b0;
            15'b01001010_0101_101: DATA = 1'b1;
            15'b01001010_0101_110: DATA = 1'b1;
            15'b01001010_0101_111: DATA = 1'b0;
            // J Row 6
            15'b01001010_0110_000: DATA = 1'b0;
            15'b01001010_0110_001: DATA = 1'b0;
            15'b01001010_0110_010: DATA = 1'b0;
            15'b01001010_0110_011: DATA = 1'b0;
            15'b01001010_0110_100: DATA = 1'b0;
            15'b01001010_0110_101: DATA = 1'b1;
            15'b01001010_0110_110: DATA = 1'b1;
            15'b01001010_0110_111: DATA = 1'b0;
            // J Row 7
            15'b01001010_0111_000: DATA = 1'b0;
            15'b01001010_0111_001: DATA = 1'b0;
            15'b01001010_0111_010: DATA = 1'b0;
            15'b01001010_0111_011: DATA = 1'b0;
            15'b01001010_0111_100: DATA = 1'b0;
            15'b01001010_0111_101: DATA = 1'b1;
            15'b01001010_0111_110: DATA = 1'b1;
            15'b01001010_0111_111: DATA = 1'b0;
            // J Row 8
            15'b01001010_1000_000: DATA = 1'b0;
            15'b01001010_1000_001: DATA = 1'b0;
            15'b01001010_1000_010: DATA = 1'b0;
            15'b01001010_1000_011: DATA = 1'b0;
            15'b01001010_1000_100: DATA = 1'b0;
            15'b01001010_1000_101: DATA = 1'b1;
            15'b01001010_1000_110: DATA = 1'b1;
            15'b01001010_1000_111: DATA = 1'b0;
            // J Row 9
            15'b01001010_1001_000: DATA = 1'b0;
            15'b01001010_1001_001: DATA = 1'b0;
            15'b01001010_1001_010: DATA = 1'b0;
            15'b01001010_1001_011: DATA = 1'b0;
            15'b01001010_1001_100: DATA = 1'b0;
            15'b01001010_1001_101: DATA = 1'b1;
            15'b01001010_1001_110: DATA = 1'b1;
            15'b01001010_1001_111: DATA = 1'b0;
            // J Row 10
            15'b01001010_1010_000: DATA = 1'b1;
            15'b01001010_1010_001: DATA = 1'b1;
            15'b01001010_1010_010: DATA = 1'b0;
            15'b01001010_1010_011: DATA = 1'b0;
            15'b01001010_1010_100: DATA = 1'b0;
            15'b01001010_1010_101: DATA = 1'b1;
            15'b01001010_1010_110: DATA = 1'b1;
            15'b01001010_1010_111: DATA = 1'b0;
            // J Row 11
            15'b01001010_1011_000: DATA = 1'b1;
            15'b01001010_1011_001: DATA = 1'b1;
            15'b01001010_1011_010: DATA = 1'b1;
            15'b01001010_1011_011: DATA = 1'b1;
            15'b01001010_1011_100: DATA = 1'b1;
            15'b01001010_1011_101: DATA = 1'b1;
            15'b01001010_1011_110: DATA = 1'b0;
            15'b01001010_1011_111: DATA = 1'b0;
            // J Row 12
            15'b01001010_1100_000: DATA = 1'b0;
            15'b01001010_1100_001: DATA = 1'b0;
            15'b01001010_1100_010: DATA = 1'b1;
            15'b01001010_1100_011: DATA = 1'b1;
            15'b01001010_1100_100: DATA = 1'b1;
            15'b01001010_1100_101: DATA = 1'b0;
            15'b01001010_1100_110: DATA = 1'b0;
            15'b01001010_1100_111: DATA = 1'b0;
            // J Row 13
            15'b01001010_1101_000: DATA = 1'b0;
            15'b01001010_1101_001: DATA = 1'b0;
            15'b01001010_1101_010: DATA = 1'b0;
            15'b01001010_1101_011: DATA = 1'b0;
            15'b01001010_1101_100: DATA = 1'b0;
            15'b01001010_1101_101: DATA = 1'b0;
            15'b01001010_1101_110: DATA = 1'b0;
            15'b01001010_1101_111: DATA = 1'b0;
            // J Row 14
            15'b01001010_1110_000: DATA = 1'b0;
            15'b01001010_1110_001: DATA = 1'b0;
            15'b01001010_1110_010: DATA = 1'b0;
            15'b01001010_1110_011: DATA = 1'b0;
            15'b01001010_1110_100: DATA = 1'b0;
            15'b01001010_1110_101: DATA = 1'b0;
            15'b01001010_1110_110: DATA = 1'b0;
            15'b01001010_1110_111: DATA = 1'b0;
            // J Row 15
            15'b01001010_1111_000: DATA = 1'b0;
            15'b01001010_1111_001: DATA = 1'b0;
            15'b01001010_1111_010: DATA = 1'b0;
            15'b01001010_1111_011: DATA = 1'b0;
            15'b01001010_1111_100: DATA = 1'b0;
            15'b01001010_1111_101: DATA = 1'b0;
            15'b01001010_1111_110: DATA = 1'b0;
            15'b01001010_1111_111: DATA = 1'b0;
            // K Row 0
            15'b01001011_0000_000: DATA = 1'b0;
            15'b01001011_0000_001: DATA = 1'b0;
            15'b01001011_0000_010: DATA = 1'b0;
            15'b01001011_0000_011: DATA = 1'b0;
            15'b01001011_0000_100: DATA = 1'b0;
            15'b01001011_0000_101: DATA = 1'b0;
            15'b01001011_0000_110: DATA = 1'b0;
            15'b01001011_0000_111: DATA = 1'b0;
            // K Row 1
            15'b01001011_0001_000: DATA = 1'b0;
            15'b01001011_0001_001: DATA = 1'b0;
            15'b01001011_0001_010: DATA = 1'b0;
            15'b01001011_0001_011: DATA = 1'b0;
            15'b01001011_0001_100: DATA = 1'b0;
            15'b01001011_0001_101: DATA = 1'b0;
            15'b01001011_0001_110: DATA = 1'b0;
            15'b01001011_0001_111: DATA = 1'b0;
            // K Row 2
            15'b01001011_0010_000: DATA = 1'b0;
            15'b01001011_0010_001: DATA = 1'b0;
            15'b01001011_0010_010: DATA = 1'b0;
            15'b01001011_0010_011: DATA = 1'b0;
            15'b01001011_0010_100: DATA = 1'b0;
            15'b01001011_0010_101: DATA = 1'b0;
            15'b01001011_0010_110: DATA = 1'b0;
            15'b01001011_0010_111: DATA = 1'b0;
            // K Row 3
            15'b01001011_0011_000: DATA = 1'b1;
            15'b01001011_0011_001: DATA = 1'b1;
            15'b01001011_0011_010: DATA = 1'b0;
            15'b01001011_0011_011: DATA = 1'b0;
            15'b01001011_0011_100: DATA = 1'b0;
            15'b01001011_0011_101: DATA = 1'b1;
            15'b01001011_0011_110: DATA = 1'b1;
            15'b01001011_0011_111: DATA = 1'b0;
            // K Row 4
            15'b01001011_0100_000: DATA = 1'b1;
            15'b01001011_0100_001: DATA = 1'b1;
            15'b01001011_0100_010: DATA = 1'b0;
            15'b01001011_0100_011: DATA = 1'b0;
            15'b01001011_0100_100: DATA = 1'b1;
            15'b01001011_0100_101: DATA = 1'b1;
            15'b01001011_0100_110: DATA = 1'b0;
            15'b01001011_0100_111: DATA = 1'b0;
            // K Row 5
            15'b01001011_0101_000: DATA = 1'b1;
            15'b01001011_0101_001: DATA = 1'b1;
            15'b01001011_0101_010: DATA = 1'b0;
            15'b01001011_0101_011: DATA = 1'b1;
            15'b01001011_0101_100: DATA = 1'b1;
            15'b01001011_0101_101: DATA = 1'b1;
            15'b01001011_0101_110: DATA = 1'b0;
            15'b01001011_0101_111: DATA = 1'b0;
            // K Row 6
            15'b01001011_0110_000: DATA = 1'b1;
            15'b01001011_0110_001: DATA = 1'b1;
            15'b01001011_0110_010: DATA = 1'b0;
            15'b01001011_0110_011: DATA = 1'b1;
            15'b01001011_0110_100: DATA = 1'b1;
            15'b01001011_0110_101: DATA = 1'b0;
            15'b01001011_0110_110: DATA = 1'b0;
            15'b01001011_0110_111: DATA = 1'b0;
            // K Row 7
            15'b01001011_0111_000: DATA = 1'b1;
            15'b01001011_0111_001: DATA = 1'b1;
            15'b01001011_0111_010: DATA = 1'b1;
            15'b01001011_0111_011: DATA = 1'b1;
            15'b01001011_0111_100: DATA = 1'b0;
            15'b01001011_0111_101: DATA = 1'b0;
            15'b01001011_0111_110: DATA = 1'b0;
            15'b01001011_0111_111: DATA = 1'b0;
            // K Row 8
            15'b01001011_1000_000: DATA = 1'b1;
            15'b01001011_1000_001: DATA = 1'b1;
            15'b01001011_1000_010: DATA = 1'b1;
            15'b01001011_1000_011: DATA = 1'b1;
            15'b01001011_1000_100: DATA = 1'b1;
            15'b01001011_1000_101: DATA = 1'b0;
            15'b01001011_1000_110: DATA = 1'b0;
            15'b01001011_1000_111: DATA = 1'b0;
            // K Row 9
            15'b01001011_1001_000: DATA = 1'b1;
            15'b01001011_1001_001: DATA = 1'b1;
            15'b01001011_1001_010: DATA = 1'b0;
            15'b01001011_1001_011: DATA = 1'b1;
            15'b01001011_1001_100: DATA = 1'b1;
            15'b01001011_1001_101: DATA = 1'b0;
            15'b01001011_1001_110: DATA = 1'b0;
            15'b01001011_1001_111: DATA = 1'b0;
            // K Row 10
            15'b01001011_1010_000: DATA = 1'b1;
            15'b01001011_1010_001: DATA = 1'b1;
            15'b01001011_1010_010: DATA = 1'b0;
            15'b01001011_1010_011: DATA = 1'b1;
            15'b01001011_1010_100: DATA = 1'b1;
            15'b01001011_1010_101: DATA = 1'b1;
            15'b01001011_1010_110: DATA = 1'b0;
            15'b01001011_1010_111: DATA = 1'b0;
            // K Row 11
            15'b01001011_1011_000: DATA = 1'b1;
            15'b01001011_1011_001: DATA = 1'b1;
            15'b01001011_1011_010: DATA = 1'b0;
            15'b01001011_1011_011: DATA = 1'b0;
            15'b01001011_1011_100: DATA = 1'b1;
            15'b01001011_1011_101: DATA = 1'b1;
            15'b01001011_1011_110: DATA = 1'b0;
            15'b01001011_1011_111: DATA = 1'b0;
            // K Row 12
            15'b01001011_1100_000: DATA = 1'b1;
            15'b01001011_1100_001: DATA = 1'b1;
            15'b01001011_1100_010: DATA = 1'b0;
            15'b01001011_1100_011: DATA = 1'b0;
            15'b01001011_1100_100: DATA = 1'b0;
            15'b01001011_1100_101: DATA = 1'b1;
            15'b01001011_1100_110: DATA = 1'b1;
            15'b01001011_1100_111: DATA = 1'b0;
            // K Row 13
            15'b01001011_1101_000: DATA = 1'b0;
            15'b01001011_1101_001: DATA = 1'b0;
            15'b01001011_1101_010: DATA = 1'b0;
            15'b01001011_1101_011: DATA = 1'b0;
            15'b01001011_1101_100: DATA = 1'b0;
            15'b01001011_1101_101: DATA = 1'b0;
            15'b01001011_1101_110: DATA = 1'b0;
            15'b01001011_1101_111: DATA = 1'b0;
            // K Row 14
            15'b01001011_1110_000: DATA = 1'b0;
            15'b01001011_1110_001: DATA = 1'b0;
            15'b01001011_1110_010: DATA = 1'b0;
            15'b01001011_1110_011: DATA = 1'b0;
            15'b01001011_1110_100: DATA = 1'b0;
            15'b01001011_1110_101: DATA = 1'b0;
            15'b01001011_1110_110: DATA = 1'b0;
            15'b01001011_1110_111: DATA = 1'b0;
            // K Row 15
            15'b01001011_1111_000: DATA = 1'b0;
            15'b01001011_1111_001: DATA = 1'b0;
            15'b01001011_1111_010: DATA = 1'b0;
            15'b01001011_1111_011: DATA = 1'b0;
            15'b01001011_1111_100: DATA = 1'b0;
            15'b01001011_1111_101: DATA = 1'b0;
            15'b01001011_1111_110: DATA = 1'b0;
            15'b01001011_1111_111: DATA = 1'b0;
            // L Row 0
            15'b01001100_0000_000: DATA = 1'b0;
            15'b01001100_0000_001: DATA = 1'b0;
            15'b01001100_0000_010: DATA = 1'b0;
            15'b01001100_0000_011: DATA = 1'b0;
            15'b01001100_0000_100: DATA = 1'b0;
            15'b01001100_0000_101: DATA = 1'b0;
            15'b01001100_0000_110: DATA = 1'b0;
            15'b01001100_0000_111: DATA = 1'b0;
            // L Row 1
            15'b01001100_0001_000: DATA = 1'b0;
            15'b01001100_0001_001: DATA = 1'b0;
            15'b01001100_0001_010: DATA = 1'b0;
            15'b01001100_0001_011: DATA = 1'b0;
            15'b01001100_0001_100: DATA = 1'b0;
            15'b01001100_0001_101: DATA = 1'b0;
            15'b01001100_0001_110: DATA = 1'b0;
            15'b01001100_0001_111: DATA = 1'b0;
            // L Row 2
            15'b01001100_0010_000: DATA = 1'b0;
            15'b01001100_0010_001: DATA = 1'b0;
            15'b01001100_0010_010: DATA = 1'b0;
            15'b01001100_0010_011: DATA = 1'b0;
            15'b01001100_0010_100: DATA = 1'b0;
            15'b01001100_0010_101: DATA = 1'b0;
            15'b01001100_0010_110: DATA = 1'b0;
            15'b01001100_0010_111: DATA = 1'b0;
            // L Row 3
            15'b01001100_0011_000: DATA = 1'b1;
            15'b01001100_0011_001: DATA = 1'b1;
            15'b01001100_0011_010: DATA = 1'b0;
            15'b01001100_0011_011: DATA = 1'b0;
            15'b01001100_0011_100: DATA = 1'b0;
            15'b01001100_0011_101: DATA = 1'b0;
            15'b01001100_0011_110: DATA = 1'b0;
            15'b01001100_0011_111: DATA = 1'b0;
            // L Row 4
            15'b01001100_0100_000: DATA = 1'b1;
            15'b01001100_0100_001: DATA = 1'b1;
            15'b01001100_0100_010: DATA = 1'b0;
            15'b01001100_0100_011: DATA = 1'b0;
            15'b01001100_0100_100: DATA = 1'b0;
            15'b01001100_0100_101: DATA = 1'b0;
            15'b01001100_0100_110: DATA = 1'b0;
            15'b01001100_0100_111: DATA = 1'b0;
            // L Row 5
            15'b01001100_0101_000: DATA = 1'b1;
            15'b01001100_0101_001: DATA = 1'b1;
            15'b01001100_0101_010: DATA = 1'b0;
            15'b01001100_0101_011: DATA = 1'b0;
            15'b01001100_0101_100: DATA = 1'b0;
            15'b01001100_0101_101: DATA = 1'b0;
            15'b01001100_0101_110: DATA = 1'b0;
            15'b01001100_0101_111: DATA = 1'b0;
            // L Row 6
            15'b01001100_0110_000: DATA = 1'b1;
            15'b01001100_0110_001: DATA = 1'b1;
            15'b01001100_0110_010: DATA = 1'b0;
            15'b01001100_0110_011: DATA = 1'b0;
            15'b01001100_0110_100: DATA = 1'b0;
            15'b01001100_0110_101: DATA = 1'b0;
            15'b01001100_0110_110: DATA = 1'b0;
            15'b01001100_0110_111: DATA = 1'b0;
            // L Row 7
            15'b01001100_0111_000: DATA = 1'b1;
            15'b01001100_0111_001: DATA = 1'b1;
            15'b01001100_0111_010: DATA = 1'b0;
            15'b01001100_0111_011: DATA = 1'b0;
            15'b01001100_0111_100: DATA = 1'b0;
            15'b01001100_0111_101: DATA = 1'b0;
            15'b01001100_0111_110: DATA = 1'b0;
            15'b01001100_0111_111: DATA = 1'b0;
            // L Row 8
            15'b01001100_1000_000: DATA = 1'b1;
            15'b01001100_1000_001: DATA = 1'b1;
            15'b01001100_1000_010: DATA = 1'b0;
            15'b01001100_1000_011: DATA = 1'b0;
            15'b01001100_1000_100: DATA = 1'b0;
            15'b01001100_1000_101: DATA = 1'b0;
            15'b01001100_1000_110: DATA = 1'b0;
            15'b01001100_1000_111: DATA = 1'b0;
            // L Row 9
            15'b01001100_1001_000: DATA = 1'b1;
            15'b01001100_1001_001: DATA = 1'b1;
            15'b01001100_1001_010: DATA = 1'b0;
            15'b01001100_1001_011: DATA = 1'b0;
            15'b01001100_1001_100: DATA = 1'b0;
            15'b01001100_1001_101: DATA = 1'b0;
            15'b01001100_1001_110: DATA = 1'b0;
            15'b01001100_1001_111: DATA = 1'b0;
            // L Row 10
            15'b01001100_1010_000: DATA = 1'b1;
            15'b01001100_1010_001: DATA = 1'b1;
            15'b01001100_1010_010: DATA = 1'b0;
            15'b01001100_1010_011: DATA = 1'b0;
            15'b01001100_1010_100: DATA = 1'b0;
            15'b01001100_1010_101: DATA = 1'b0;
            15'b01001100_1010_110: DATA = 1'b0;
            15'b01001100_1010_111: DATA = 1'b0;
            // L Row 11
            15'b01001100_1011_000: DATA = 1'b1;
            15'b01001100_1011_001: DATA = 1'b1;
            15'b01001100_1011_010: DATA = 1'b1;
            15'b01001100_1011_011: DATA = 1'b1;
            15'b01001100_1011_100: DATA = 1'b1;
            15'b01001100_1011_101: DATA = 1'b1;
            15'b01001100_1011_110: DATA = 1'b1;
            15'b01001100_1011_111: DATA = 1'b0;
            // L Row 12
            15'b01001100_1100_000: DATA = 1'b1;
            15'b01001100_1100_001: DATA = 1'b1;
            15'b01001100_1100_010: DATA = 1'b1;
            15'b01001100_1100_011: DATA = 1'b1;
            15'b01001100_1100_100: DATA = 1'b1;
            15'b01001100_1100_101: DATA = 1'b1;
            15'b01001100_1100_110: DATA = 1'b1;
            15'b01001100_1100_111: DATA = 1'b0;
            // L Row 13
            15'b01001100_1101_000: DATA = 1'b0;
            15'b01001100_1101_001: DATA = 1'b0;
            15'b01001100_1101_010: DATA = 1'b0;
            15'b01001100_1101_011: DATA = 1'b0;
            15'b01001100_1101_100: DATA = 1'b0;
            15'b01001100_1101_101: DATA = 1'b0;
            15'b01001100_1101_110: DATA = 1'b0;
            15'b01001100_1101_111: DATA = 1'b0;
            // L Row 14
            15'b01001100_1110_000: DATA = 1'b0;
            15'b01001100_1110_001: DATA = 1'b0;
            15'b01001100_1110_010: DATA = 1'b0;
            15'b01001100_1110_011: DATA = 1'b0;
            15'b01001100_1110_100: DATA = 1'b0;
            15'b01001100_1110_101: DATA = 1'b0;
            15'b01001100_1110_110: DATA = 1'b0;
            15'b01001100_1110_111: DATA = 1'b0;
            // L Row 15
            15'b01001100_1111_000: DATA = 1'b0;
            15'b01001100_1111_001: DATA = 1'b0;
            15'b01001100_1111_010: DATA = 1'b0;
            15'b01001100_1111_011: DATA = 1'b0;
            15'b01001100_1111_100: DATA = 1'b0;
            15'b01001100_1111_101: DATA = 1'b0;
            15'b01001100_1111_110: DATA = 1'b0;
            15'b01001100_1111_111: DATA = 1'b0;
            // M Row 0
            15'b01001101_0000_000: DATA = 1'b0;
            15'b01001101_0000_001: DATA = 1'b0;
            15'b01001101_0000_010: DATA = 1'b0;
            15'b01001101_0000_011: DATA = 1'b0;
            15'b01001101_0000_100: DATA = 1'b0;
            15'b01001101_0000_101: DATA = 1'b0;
            15'b01001101_0000_110: DATA = 1'b0;
            15'b01001101_0000_111: DATA = 1'b0;
            // M Row 1
            15'b01001101_0001_000: DATA = 1'b0;
            15'b01001101_0001_001: DATA = 1'b0;
            15'b01001101_0001_010: DATA = 1'b0;
            15'b01001101_0001_011: DATA = 1'b0;
            15'b01001101_0001_100: DATA = 1'b0;
            15'b01001101_0001_101: DATA = 1'b0;
            15'b01001101_0001_110: DATA = 1'b0;
            15'b01001101_0001_111: DATA = 1'b0;
            // M Row 2
            15'b01001101_0010_000: DATA = 1'b0;
            15'b01001101_0010_001: DATA = 1'b0;
            15'b01001101_0010_010: DATA = 1'b0;
            15'b01001101_0010_011: DATA = 1'b0;
            15'b01001101_0010_100: DATA = 1'b0;
            15'b01001101_0010_101: DATA = 1'b0;
            15'b01001101_0010_110: DATA = 1'b0;
            15'b01001101_0010_111: DATA = 1'b0;
            // M Row 3
            15'b01001101_0011_000: DATA = 1'b1;
            15'b01001101_0011_001: DATA = 1'b1;
            15'b01001101_0011_010: DATA = 1'b0;
            15'b01001101_0011_011: DATA = 1'b0;
            15'b01001101_0011_100: DATA = 1'b0;
            15'b01001101_0011_101: DATA = 1'b1;
            15'b01001101_0011_110: DATA = 1'b1;
            15'b01001101_0011_111: DATA = 1'b0;
            // M Row 4
            15'b01001101_0100_000: DATA = 1'b1;
            15'b01001101_0100_001: DATA = 1'b1;
            15'b01001101_0100_010: DATA = 1'b1;
            15'b01001101_0100_011: DATA = 1'b0;
            15'b01001101_0100_100: DATA = 1'b1;
            15'b01001101_0100_101: DATA = 1'b1;
            15'b01001101_0100_110: DATA = 1'b1;
            15'b01001101_0100_111: DATA = 1'b0;
            // M Row 5
            15'b01001101_0101_000: DATA = 1'b1;
            15'b01001101_0101_001: DATA = 1'b1;
            15'b01001101_0101_010: DATA = 1'b1;
            15'b01001101_0101_011: DATA = 1'b1;
            15'b01001101_0101_100: DATA = 1'b1;
            15'b01001101_0101_101: DATA = 1'b0;
            15'b01001101_0101_110: DATA = 1'b1;
            15'b01001101_0101_111: DATA = 1'b0;
            // M Row 6
            15'b01001101_0110_000: DATA = 1'b1;
            15'b01001101_0110_001: DATA = 1'b1;
            15'b01001101_0110_010: DATA = 1'b0;
            15'b01001101_0110_011: DATA = 1'b1;
            15'b01001101_0110_100: DATA = 1'b1;
            15'b01001101_0110_101: DATA = 1'b0;
            15'b01001101_0110_110: DATA = 1'b1;
            15'b01001101_0110_111: DATA = 1'b0;
            // M Row 7
            15'b01001101_0111_000: DATA = 1'b1;
            15'b01001101_0111_001: DATA = 1'b1;
            15'b01001101_0111_010: DATA = 1'b0;
            15'b01001101_0111_011: DATA = 1'b1;
            15'b01001101_0111_100: DATA = 1'b0;
            15'b01001101_0111_101: DATA = 1'b0;
            15'b01001101_0111_110: DATA = 1'b1;
            15'b01001101_0111_111: DATA = 1'b0;
            // M Row 8
            15'b01001101_1000_000: DATA = 1'b1;
            15'b01001101_1000_001: DATA = 1'b1;
            15'b01001101_1000_010: DATA = 1'b0;
            15'b01001101_1000_011: DATA = 1'b0;
            15'b01001101_1000_100: DATA = 1'b0;
            15'b01001101_1000_101: DATA = 1'b0;
            15'b01001101_1000_110: DATA = 1'b1;
            15'b01001101_1000_111: DATA = 1'b0;
            // M Row 9
            15'b01001101_1001_000: DATA = 1'b1;
            15'b01001101_1001_001: DATA = 1'b1;
            15'b01001101_1001_010: DATA = 1'b0;
            15'b01001101_1001_011: DATA = 1'b0;
            15'b01001101_1001_100: DATA = 1'b0;
            15'b01001101_1001_101: DATA = 1'b0;
            15'b01001101_1001_110: DATA = 1'b1;
            15'b01001101_1001_111: DATA = 1'b0;
            // M Row 10
            15'b01001101_1010_000: DATA = 1'b1;
            15'b01001101_1010_001: DATA = 1'b1;
            15'b01001101_1010_010: DATA = 1'b0;
            15'b01001101_1010_011: DATA = 1'b0;
            15'b01001101_1010_100: DATA = 1'b0;
            15'b01001101_1010_101: DATA = 1'b0;
            15'b01001101_1010_110: DATA = 1'b1;
            15'b01001101_1010_111: DATA = 1'b0;
            // M Row 11
            15'b01001101_1011_000: DATA = 1'b1;
            15'b01001101_1011_001: DATA = 1'b1;
            15'b01001101_1011_010: DATA = 1'b0;
            15'b01001101_1011_011: DATA = 1'b0;
            15'b01001101_1011_100: DATA = 1'b0;
            15'b01001101_1011_101: DATA = 1'b0;
            15'b01001101_1011_110: DATA = 1'b1;
            15'b01001101_1011_111: DATA = 1'b0;
            // M Row 12
            15'b01001101_1100_000: DATA = 1'b1;
            15'b01001101_1100_001: DATA = 1'b1;
            15'b01001101_1100_010: DATA = 1'b0;
            15'b01001101_1100_011: DATA = 1'b0;
            15'b01001101_1100_100: DATA = 1'b0;
            15'b01001101_1100_101: DATA = 1'b0;
            15'b01001101_1100_110: DATA = 1'b1;
            15'b01001101_1100_111: DATA = 1'b0;
            // M Row 13
            15'b01001101_1101_000: DATA = 1'b0;
            15'b01001101_1101_001: DATA = 1'b0;
            15'b01001101_1101_010: DATA = 1'b0;
            15'b01001101_1101_011: DATA = 1'b0;
            15'b01001101_1101_100: DATA = 1'b0;
            15'b01001101_1101_101: DATA = 1'b0;
            15'b01001101_1101_110: DATA = 1'b0;
            15'b01001101_1101_111: DATA = 1'b0;
            // M Row 14
            15'b01001101_1110_000: DATA = 1'b0;
            15'b01001101_1110_001: DATA = 1'b0;
            15'b01001101_1110_010: DATA = 1'b0;
            15'b01001101_1110_011: DATA = 1'b0;
            15'b01001101_1110_100: DATA = 1'b0;
            15'b01001101_1110_101: DATA = 1'b0;
            15'b01001101_1110_110: DATA = 1'b0;
            15'b01001101_1110_111: DATA = 1'b0;
            // M Row 15
            15'b01001101_1111_000: DATA = 1'b0;
            15'b01001101_1111_001: DATA = 1'b0;
            15'b01001101_1111_010: DATA = 1'b0;
            15'b01001101_1111_011: DATA = 1'b0;
            15'b01001101_1111_100: DATA = 1'b0;
            15'b01001101_1111_101: DATA = 1'b0;
            15'b01001101_1111_110: DATA = 1'b0;
            15'b01001101_1111_111: DATA = 1'b0;
            // N Row 0
            15'b01001110_0000_000: DATA = 1'b0;
            15'b01001110_0000_001: DATA = 1'b0;
            15'b01001110_0000_010: DATA = 1'b0;
            15'b01001110_0000_011: DATA = 1'b0;
            15'b01001110_0000_100: DATA = 1'b0;
            15'b01001110_0000_101: DATA = 1'b0;
            15'b01001110_0000_110: DATA = 1'b0;
            15'b01001110_0000_111: DATA = 1'b0;
            // N Row 1
            15'b01001110_0001_000: DATA = 1'b0;
            15'b01001110_0001_001: DATA = 1'b0;
            15'b01001110_0001_010: DATA = 1'b0;
            15'b01001110_0001_011: DATA = 1'b0;
            15'b01001110_0001_100: DATA = 1'b0;
            15'b01001110_0001_101: DATA = 1'b0;
            15'b01001110_0001_110: DATA = 1'b0;
            15'b01001110_0001_111: DATA = 1'b0;
            // N Row 2
            15'b01001110_0010_000: DATA = 1'b0;
            15'b01001110_0010_001: DATA = 1'b0;
            15'b01001110_0010_010: DATA = 1'b0;
            15'b01001110_0010_011: DATA = 1'b0;
            15'b01001110_0010_100: DATA = 1'b0;
            15'b01001110_0010_101: DATA = 1'b0;
            15'b01001110_0010_110: DATA = 1'b0;
            15'b01001110_0010_111: DATA = 1'b0;
            // N Row 3
            15'b01001110_0011_000: DATA = 1'b1;
            15'b01001110_0011_001: DATA = 1'b1;
            15'b01001110_0011_010: DATA = 1'b1;
            15'b01001110_0011_011: DATA = 1'b0;
            15'b01001110_0011_100: DATA = 1'b0;
            15'b01001110_0011_101: DATA = 1'b0;
            15'b01001110_0011_110: DATA = 1'b1;
            15'b01001110_0011_111: DATA = 1'b0;
            // N Row 4
            15'b01001110_0100_000: DATA = 1'b1;
            15'b01001110_0100_001: DATA = 1'b1;
            15'b01001110_0100_010: DATA = 1'b1;
            15'b01001110_0100_011: DATA = 1'b0;
            15'b01001110_0100_100: DATA = 1'b0;
            15'b01001110_0100_101: DATA = 1'b0;
            15'b01001110_0100_110: DATA = 1'b1;
            15'b01001110_0100_111: DATA = 1'b0;
            // N Row 5
            15'b01001110_0101_000: DATA = 1'b1;
            15'b01001110_0101_001: DATA = 1'b1;
            15'b01001110_0101_010: DATA = 1'b1;
            15'b01001110_0101_011: DATA = 1'b1;
            15'b01001110_0101_100: DATA = 1'b0;
            15'b01001110_0101_101: DATA = 1'b0;
            15'b01001110_0101_110: DATA = 1'b1;
            15'b01001110_0101_111: DATA = 1'b0;
            // N Row 6
            15'b01001110_0110_000: DATA = 1'b1;
            15'b01001110_0110_001: DATA = 1'b1;
            15'b01001110_0110_010: DATA = 1'b0;
            15'b01001110_0110_011: DATA = 1'b1;
            15'b01001110_0110_100: DATA = 1'b1;
            15'b01001110_0110_101: DATA = 1'b0;
            15'b01001110_0110_110: DATA = 1'b1;
            15'b01001110_0110_111: DATA = 1'b0;
            // N Row 7
            15'b01001110_0111_000: DATA = 1'b1;
            15'b01001110_0111_001: DATA = 1'b1;
            15'b01001110_0111_010: DATA = 1'b0;
            15'b01001110_0111_011: DATA = 1'b1;
            15'b01001110_0111_100: DATA = 1'b1;
            15'b01001110_0111_101: DATA = 1'b0;
            15'b01001110_0111_110: DATA = 1'b1;
            15'b01001110_0111_111: DATA = 1'b0;
            // N Row 8
            15'b01001110_1000_000: DATA = 1'b1;
            15'b01001110_1000_001: DATA = 1'b1;
            15'b01001110_1000_010: DATA = 1'b0;
            15'b01001110_1000_011: DATA = 1'b1;
            15'b01001110_1000_100: DATA = 1'b1;
            15'b01001110_1000_101: DATA = 1'b0;
            15'b01001110_1000_110: DATA = 1'b1;
            15'b01001110_1000_111: DATA = 1'b0;
            // N Row 9
            15'b01001110_1001_000: DATA = 1'b1;
            15'b01001110_1001_001: DATA = 1'b1;
            15'b01001110_1001_010: DATA = 1'b0;
            15'b01001110_1001_011: DATA = 1'b0;
            15'b01001110_1001_100: DATA = 1'b1;
            15'b01001110_1001_101: DATA = 1'b0;
            15'b01001110_1001_110: DATA = 1'b1;
            15'b01001110_1001_111: DATA = 1'b0;
            // N Row 10
            15'b01001110_1010_000: DATA = 1'b1;
            15'b01001110_1010_001: DATA = 1'b1;
            15'b01001110_1010_010: DATA = 1'b0;
            15'b01001110_1010_011: DATA = 1'b0;
            15'b01001110_1010_100: DATA = 1'b1;
            15'b01001110_1010_101: DATA = 1'b1;
            15'b01001110_1010_110: DATA = 1'b1;
            15'b01001110_1010_111: DATA = 1'b0;
            // N Row 11
            15'b01001110_1011_000: DATA = 1'b1;
            15'b01001110_1011_001: DATA = 1'b1;
            15'b01001110_1011_010: DATA = 1'b0;
            15'b01001110_1011_011: DATA = 1'b0;
            15'b01001110_1011_100: DATA = 1'b0;
            15'b01001110_1011_101: DATA = 1'b1;
            15'b01001110_1011_110: DATA = 1'b1;
            15'b01001110_1011_111: DATA = 1'b0;
            // N Row 12
            15'b01001110_1100_000: DATA = 1'b1;
            15'b01001110_1100_001: DATA = 1'b1;
            15'b01001110_1100_010: DATA = 1'b0;
            15'b01001110_1100_011: DATA = 1'b0;
            15'b01001110_1100_100: DATA = 1'b0;
            15'b01001110_1100_101: DATA = 1'b1;
            15'b01001110_1100_110: DATA = 1'b1;
            15'b01001110_1100_111: DATA = 1'b0;
            // N Row 13
            15'b01001110_1101_000: DATA = 1'b0;
            15'b01001110_1101_001: DATA = 1'b0;
            15'b01001110_1101_010: DATA = 1'b0;
            15'b01001110_1101_011: DATA = 1'b0;
            15'b01001110_1101_100: DATA = 1'b0;
            15'b01001110_1101_101: DATA = 1'b0;
            15'b01001110_1101_110: DATA = 1'b0;
            15'b01001110_1101_111: DATA = 1'b0;
            // N Row 14
            15'b01001110_1110_000: DATA = 1'b0;
            15'b01001110_1110_001: DATA = 1'b0;
            15'b01001110_1110_010: DATA = 1'b0;
            15'b01001110_1110_011: DATA = 1'b0;
            15'b01001110_1110_100: DATA = 1'b0;
            15'b01001110_1110_101: DATA = 1'b0;
            15'b01001110_1110_110: DATA = 1'b0;
            15'b01001110_1110_111: DATA = 1'b0;
            // N Row 15
            15'b01001110_1111_000: DATA = 1'b0;
            15'b01001110_1111_001: DATA = 1'b0;
            15'b01001110_1111_010: DATA = 1'b0;
            15'b01001110_1111_011: DATA = 1'b0;
            15'b01001110_1111_100: DATA = 1'b0;
            15'b01001110_1111_101: DATA = 1'b0;
            15'b01001110_1111_110: DATA = 1'b0;
            15'b01001110_1111_111: DATA = 1'b0;
            // O Row 0
            15'b01001111_0000_000: DATA = 1'b0;
            15'b01001111_0000_001: DATA = 1'b0;
            15'b01001111_0000_010: DATA = 1'b0;
            15'b01001111_0000_011: DATA = 1'b0;
            15'b01001111_0000_100: DATA = 1'b0;
            15'b01001111_0000_101: DATA = 1'b0;
            15'b01001111_0000_110: DATA = 1'b0;
            15'b01001111_0000_111: DATA = 1'b0;
            // O Row 1
            15'b01001111_0001_000: DATA = 1'b0;
            15'b01001111_0001_001: DATA = 1'b0;
            15'b01001111_0001_010: DATA = 1'b0;
            15'b01001111_0001_011: DATA = 1'b0;
            15'b01001111_0001_100: DATA = 1'b0;
            15'b01001111_0001_101: DATA = 1'b0;
            15'b01001111_0001_110: DATA = 1'b0;
            15'b01001111_0001_111: DATA = 1'b0;
            // O Row 2
            15'b01001111_0010_000: DATA = 1'b0;
            15'b01001111_0010_001: DATA = 1'b0;
            15'b01001111_0010_010: DATA = 1'b0;
            15'b01001111_0010_011: DATA = 1'b0;
            15'b01001111_0010_100: DATA = 1'b0;
            15'b01001111_0010_101: DATA = 1'b0;
            15'b01001111_0010_110: DATA = 1'b0;
            15'b01001111_0010_111: DATA = 1'b0;
            // O Row 3
            15'b01001111_0011_000: DATA = 1'b0;
            15'b01001111_0011_001: DATA = 1'b0;
            15'b01001111_0011_010: DATA = 1'b1;
            15'b01001111_0011_011: DATA = 1'b1;
            15'b01001111_0011_100: DATA = 1'b1;
            15'b01001111_0011_101: DATA = 1'b0;
            15'b01001111_0011_110: DATA = 1'b0;
            15'b01001111_0011_111: DATA = 1'b0;
            // O Row 4
            15'b01001111_0100_000: DATA = 1'b0;
            15'b01001111_0100_001: DATA = 1'b1;
            15'b01001111_0100_010: DATA = 1'b1;
            15'b01001111_0100_011: DATA = 1'b1;
            15'b01001111_0100_100: DATA = 1'b1;
            15'b01001111_0100_101: DATA = 1'b1;
            15'b01001111_0100_110: DATA = 1'b0;
            15'b01001111_0100_111: DATA = 1'b0;
            // O Row 5
            15'b01001111_0101_000: DATA = 1'b1;
            15'b01001111_0101_001: DATA = 1'b1;
            15'b01001111_0101_010: DATA = 1'b0;
            15'b01001111_0101_011: DATA = 1'b0;
            15'b01001111_0101_100: DATA = 1'b0;
            15'b01001111_0101_101: DATA = 1'b1;
            15'b01001111_0101_110: DATA = 1'b1;
            15'b01001111_0101_111: DATA = 1'b0;
            // O Row 6
            15'b01001111_0110_000: DATA = 1'b1;
            15'b01001111_0110_001: DATA = 1'b1;
            15'b01001111_0110_010: DATA = 1'b0;
            15'b01001111_0110_011: DATA = 1'b0;
            15'b01001111_0110_100: DATA = 1'b0;
            15'b01001111_0110_101: DATA = 1'b1;
            15'b01001111_0110_110: DATA = 1'b1;
            15'b01001111_0110_111: DATA = 1'b0;
            // O Row 7
            15'b01001111_0111_000: DATA = 1'b1;
            15'b01001111_0111_001: DATA = 1'b1;
            15'b01001111_0111_010: DATA = 1'b0;
            15'b01001111_0111_011: DATA = 1'b0;
            15'b01001111_0111_100: DATA = 1'b0;
            15'b01001111_0111_101: DATA = 1'b1;
            15'b01001111_0111_110: DATA = 1'b1;
            15'b01001111_0111_111: DATA = 1'b0;
            // O Row 8
            15'b01001111_1000_000: DATA = 1'b1;
            15'b01001111_1000_001: DATA = 1'b1;
            15'b01001111_1000_010: DATA = 1'b0;
            15'b01001111_1000_011: DATA = 1'b0;
            15'b01001111_1000_100: DATA = 1'b0;
            15'b01001111_1000_101: DATA = 1'b1;
            15'b01001111_1000_110: DATA = 1'b1;
            15'b01001111_1000_111: DATA = 1'b0;
            // O Row 9
            15'b01001111_1001_000: DATA = 1'b1;
            15'b01001111_1001_001: DATA = 1'b1;
            15'b01001111_1001_010: DATA = 1'b0;
            15'b01001111_1001_011: DATA = 1'b0;
            15'b01001111_1001_100: DATA = 1'b0;
            15'b01001111_1001_101: DATA = 1'b1;
            15'b01001111_1001_110: DATA = 1'b1;
            15'b01001111_1001_111: DATA = 1'b0;
            // O Row 10
            15'b01001111_1010_000: DATA = 1'b1;
            15'b01001111_1010_001: DATA = 1'b1;
            15'b01001111_1010_010: DATA = 1'b0;
            15'b01001111_1010_011: DATA = 1'b0;
            15'b01001111_1010_100: DATA = 1'b0;
            15'b01001111_1010_101: DATA = 1'b1;
            15'b01001111_1010_110: DATA = 1'b1;
            15'b01001111_1010_111: DATA = 1'b0;
            // O Row 11
            15'b01001111_1011_000: DATA = 1'b0;
            15'b01001111_1011_001: DATA = 1'b1;
            15'b01001111_1011_010: DATA = 1'b1;
            15'b01001111_1011_011: DATA = 1'b1;
            15'b01001111_1011_100: DATA = 1'b1;
            15'b01001111_1011_101: DATA = 1'b1;
            15'b01001111_1011_110: DATA = 1'b0;
            15'b01001111_1011_111: DATA = 1'b0;
            // O Row 12
            15'b01001111_1100_000: DATA = 1'b0;
            15'b01001111_1100_001: DATA = 1'b0;
            15'b01001111_1100_010: DATA = 1'b1;
            15'b01001111_1100_011: DATA = 1'b1;
            15'b01001111_1100_100: DATA = 1'b1;
            15'b01001111_1100_101: DATA = 1'b0;
            15'b01001111_1100_110: DATA = 1'b0;
            15'b01001111_1100_111: DATA = 1'b0;
            // O Row 13
            15'b01001111_1101_000: DATA = 1'b0;
            15'b01001111_1101_001: DATA = 1'b0;
            15'b01001111_1101_010: DATA = 1'b0;
            15'b01001111_1101_011: DATA = 1'b0;
            15'b01001111_1101_100: DATA = 1'b0;
            15'b01001111_1101_101: DATA = 1'b0;
            15'b01001111_1101_110: DATA = 1'b0;
            15'b01001111_1101_111: DATA = 1'b0;
            // O Row 14
            15'b01001111_1110_000: DATA = 1'b0;
            15'b01001111_1110_001: DATA = 1'b0;
            15'b01001111_1110_010: DATA = 1'b0;
            15'b01001111_1110_011: DATA = 1'b0;
            15'b01001111_1110_100: DATA = 1'b0;
            15'b01001111_1110_101: DATA = 1'b0;
            15'b01001111_1110_110: DATA = 1'b0;
            15'b01001111_1110_111: DATA = 1'b0;
            // O Row 15
            15'b01001111_1111_000: DATA = 1'b0;
            15'b01001111_1111_001: DATA = 1'b0;
            15'b01001111_1111_010: DATA = 1'b0;
            15'b01001111_1111_011: DATA = 1'b0;
            15'b01001111_1111_100: DATA = 1'b0;
            15'b01001111_1111_101: DATA = 1'b0;
            15'b01001111_1111_110: DATA = 1'b0;
            15'b01001111_1111_111: DATA = 1'b0;
            // P Row 0
            15'b01010000_0000_000: DATA = 1'b0;
            15'b01010000_0000_001: DATA = 1'b0;
            15'b01010000_0000_010: DATA = 1'b0;
            15'b01010000_0000_011: DATA = 1'b0;
            15'b01010000_0000_100: DATA = 1'b0;
            15'b01010000_0000_101: DATA = 1'b0;
            15'b01010000_0000_110: DATA = 1'b0;
            15'b01010000_0000_111: DATA = 1'b0;
            // P Row 1
            15'b01010000_0001_000: DATA = 1'b0;
            15'b01010000_0001_001: DATA = 1'b0;
            15'b01010000_0001_010: DATA = 1'b0;
            15'b01010000_0001_011: DATA = 1'b0;
            15'b01010000_0001_100: DATA = 1'b0;
            15'b01010000_0001_101: DATA = 1'b0;
            15'b01010000_0001_110: DATA = 1'b0;
            15'b01010000_0001_111: DATA = 1'b0;
            // P Row 2
            15'b01010000_0010_000: DATA = 1'b0;
            15'b01010000_0010_001: DATA = 1'b0;
            15'b01010000_0010_010: DATA = 1'b0;
            15'b01010000_0010_011: DATA = 1'b0;
            15'b01010000_0010_100: DATA = 1'b0;
            15'b01010000_0010_101: DATA = 1'b0;
            15'b01010000_0010_110: DATA = 1'b0;
            15'b01010000_0010_111: DATA = 1'b0;
            // P Row 3
            15'b01010000_0011_000: DATA = 1'b1;
            15'b01010000_0011_001: DATA = 1'b1;
            15'b01010000_0011_010: DATA = 1'b1;
            15'b01010000_0011_011: DATA = 1'b1;
            15'b01010000_0011_100: DATA = 1'b1;
            15'b01010000_0011_101: DATA = 1'b0;
            15'b01010000_0011_110: DATA = 1'b0;
            15'b01010000_0011_111: DATA = 1'b0;
            // P Row 4
            15'b01010000_0100_000: DATA = 1'b1;
            15'b01010000_0100_001: DATA = 1'b1;
            15'b01010000_0100_010: DATA = 1'b1;
            15'b01010000_0100_011: DATA = 1'b1;
            15'b01010000_0100_100: DATA = 1'b1;
            15'b01010000_0100_101: DATA = 1'b1;
            15'b01010000_0100_110: DATA = 1'b0;
            15'b01010000_0100_111: DATA = 1'b0;
            // P Row 5
            15'b01010000_0101_000: DATA = 1'b1;
            15'b01010000_0101_001: DATA = 1'b1;
            15'b01010000_0101_010: DATA = 1'b0;
            15'b01010000_0101_011: DATA = 1'b0;
            15'b01010000_0101_100: DATA = 1'b0;
            15'b01010000_0101_101: DATA = 1'b1;
            15'b01010000_0101_110: DATA = 1'b1;
            15'b01010000_0101_111: DATA = 1'b0;
            // P Row 6
            15'b01010000_0110_000: DATA = 1'b1;
            15'b01010000_0110_001: DATA = 1'b1;
            15'b01010000_0110_010: DATA = 1'b0;
            15'b01010000_0110_011: DATA = 1'b0;
            15'b01010000_0110_100: DATA = 1'b0;
            15'b01010000_0110_101: DATA = 1'b1;
            15'b01010000_0110_110: DATA = 1'b1;
            15'b01010000_0110_111: DATA = 1'b0;
            // P Row 7
            15'b01010000_0111_000: DATA = 1'b1;
            15'b01010000_0111_001: DATA = 1'b1;
            15'b01010000_0111_010: DATA = 1'b1;
            15'b01010000_0111_011: DATA = 1'b1;
            15'b01010000_0111_100: DATA = 1'b1;
            15'b01010000_0111_101: DATA = 1'b1;
            15'b01010000_0111_110: DATA = 1'b0;
            15'b01010000_0111_111: DATA = 1'b0;
            // P Row 8
            15'b01010000_1000_000: DATA = 1'b1;
            15'b01010000_1000_001: DATA = 1'b1;
            15'b01010000_1000_010: DATA = 1'b1;
            15'b01010000_1000_011: DATA = 1'b1;
            15'b01010000_1000_100: DATA = 1'b1;
            15'b01010000_1000_101: DATA = 1'b0;
            15'b01010000_1000_110: DATA = 1'b0;
            15'b01010000_1000_111: DATA = 1'b0;
            // P Row 9
            15'b01010000_1001_000: DATA = 1'b1;
            15'b01010000_1001_001: DATA = 1'b1;
            15'b01010000_1001_010: DATA = 1'b0;
            15'b01010000_1001_011: DATA = 1'b0;
            15'b01010000_1001_100: DATA = 1'b0;
            15'b01010000_1001_101: DATA = 1'b0;
            15'b01010000_1001_110: DATA = 1'b0;
            15'b01010000_1001_111: DATA = 1'b0;
            // P Row 10
            15'b01010000_1010_000: DATA = 1'b1;
            15'b01010000_1010_001: DATA = 1'b1;
            15'b01010000_1010_010: DATA = 1'b0;
            15'b01010000_1010_011: DATA = 1'b0;
            15'b01010000_1010_100: DATA = 1'b0;
            15'b01010000_1010_101: DATA = 1'b0;
            15'b01010000_1010_110: DATA = 1'b0;
            15'b01010000_1010_111: DATA = 1'b0;
            // P Row 11
            15'b01010000_1011_000: DATA = 1'b1;
            15'b01010000_1011_001: DATA = 1'b1;
            15'b01010000_1011_010: DATA = 1'b0;
            15'b01010000_1011_011: DATA = 1'b0;
            15'b01010000_1011_100: DATA = 1'b0;
            15'b01010000_1011_101: DATA = 1'b0;
            15'b01010000_1011_110: DATA = 1'b0;
            15'b01010000_1011_111: DATA = 1'b0;
            // P Row 12
            15'b01010000_1100_000: DATA = 1'b1;
            15'b01010000_1100_001: DATA = 1'b1;
            15'b01010000_1100_010: DATA = 1'b0;
            15'b01010000_1100_011: DATA = 1'b0;
            15'b01010000_1100_100: DATA = 1'b0;
            15'b01010000_1100_101: DATA = 1'b0;
            15'b01010000_1100_110: DATA = 1'b0;
            15'b01010000_1100_111: DATA = 1'b0;
            // P Row 13
            15'b01010000_1101_000: DATA = 1'b0;
            15'b01010000_1101_001: DATA = 1'b0;
            15'b01010000_1101_010: DATA = 1'b0;
            15'b01010000_1101_011: DATA = 1'b0;
            15'b01010000_1101_100: DATA = 1'b0;
            15'b01010000_1101_101: DATA = 1'b0;
            15'b01010000_1101_110: DATA = 1'b0;
            15'b01010000_1101_111: DATA = 1'b0;
            // P Row 14
            15'b01010000_1110_000: DATA = 1'b0;
            15'b01010000_1110_001: DATA = 1'b0;
            15'b01010000_1110_010: DATA = 1'b0;
            15'b01010000_1110_011: DATA = 1'b0;
            15'b01010000_1110_100: DATA = 1'b0;
            15'b01010000_1110_101: DATA = 1'b0;
            15'b01010000_1110_110: DATA = 1'b0;
            15'b01010000_1110_111: DATA = 1'b0;
            // P Row 15
            15'b01010000_1111_000: DATA = 1'b0;
            15'b01010000_1111_001: DATA = 1'b0;
            15'b01010000_1111_010: DATA = 1'b0;
            15'b01010000_1111_011: DATA = 1'b0;
            15'b01010000_1111_100: DATA = 1'b0;
            15'b01010000_1111_101: DATA = 1'b0;
            15'b01010000_1111_110: DATA = 1'b0;
            15'b01010000_1111_111: DATA = 1'b0;
            // Q Row 0
            15'b01010001_0000_000: DATA = 1'b0;
            15'b01010001_0000_001: DATA = 1'b0;
            15'b01010001_0000_010: DATA = 1'b0;
            15'b01010001_0000_011: DATA = 1'b0;
            15'b01010001_0000_100: DATA = 1'b0;
            15'b01010001_0000_101: DATA = 1'b0;
            15'b01010001_0000_110: DATA = 1'b0;
            15'b01010001_0000_111: DATA = 1'b0;
            // Q Row 1
            15'b01010001_0001_000: DATA = 1'b0;
            15'b01010001_0001_001: DATA = 1'b0;
            15'b01010001_0001_010: DATA = 1'b0;
            15'b01010001_0001_011: DATA = 1'b0;
            15'b01010001_0001_100: DATA = 1'b0;
            15'b01010001_0001_101: DATA = 1'b0;
            15'b01010001_0001_110: DATA = 1'b0;
            15'b01010001_0001_111: DATA = 1'b0;
            // Q Row 2
            15'b01010001_0010_000: DATA = 1'b0;
            15'b01010001_0010_001: DATA = 1'b0;
            15'b01010001_0010_010: DATA = 1'b0;
            15'b01010001_0010_011: DATA = 1'b0;
            15'b01010001_0010_100: DATA = 1'b0;
            15'b01010001_0010_101: DATA = 1'b0;
            15'b01010001_0010_110: DATA = 1'b0;
            15'b01010001_0010_111: DATA = 1'b0;
            // Q Row 3
            15'b01010001_0011_000: DATA = 1'b0;
            15'b01010001_0011_001: DATA = 1'b0;
            15'b01010001_0011_010: DATA = 1'b1;
            15'b01010001_0011_011: DATA = 1'b1;
            15'b01010001_0011_100: DATA = 1'b1;
            15'b01010001_0011_101: DATA = 1'b0;
            15'b01010001_0011_110: DATA = 1'b0;
            15'b01010001_0011_111: DATA = 1'b0;
            // Q Row 4
            15'b01010001_0100_000: DATA = 1'b0;
            15'b01010001_0100_001: DATA = 1'b1;
            15'b01010001_0100_010: DATA = 1'b1;
            15'b01010001_0100_011: DATA = 1'b1;
            15'b01010001_0100_100: DATA = 1'b1;
            15'b01010001_0100_101: DATA = 1'b1;
            15'b01010001_0100_110: DATA = 1'b0;
            15'b01010001_0100_111: DATA = 1'b0;
            // Q Row 5
            15'b01010001_0101_000: DATA = 1'b1;
            15'b01010001_0101_001: DATA = 1'b1;
            15'b01010001_0101_010: DATA = 1'b0;
            15'b01010001_0101_011: DATA = 1'b0;
            15'b01010001_0101_100: DATA = 1'b0;
            15'b01010001_0101_101: DATA = 1'b1;
            15'b01010001_0101_110: DATA = 1'b1;
            15'b01010001_0101_111: DATA = 1'b0;
            // Q Row 6
            15'b01010001_0110_000: DATA = 1'b1;
            15'b01010001_0110_001: DATA = 1'b1;
            15'b01010001_0110_010: DATA = 1'b0;
            15'b01010001_0110_011: DATA = 1'b0;
            15'b01010001_0110_100: DATA = 1'b0;
            15'b01010001_0110_101: DATA = 1'b1;
            15'b01010001_0110_110: DATA = 1'b1;
            15'b01010001_0110_111: DATA = 1'b0;
            // Q Row 7
            15'b01010001_0111_000: DATA = 1'b1;
            15'b01010001_0111_001: DATA = 1'b1;
            15'b01010001_0111_010: DATA = 1'b0;
            15'b01010001_0111_011: DATA = 1'b0;
            15'b01010001_0111_100: DATA = 1'b0;
            15'b01010001_0111_101: DATA = 1'b1;
            15'b01010001_0111_110: DATA = 1'b1;
            15'b01010001_0111_111: DATA = 1'b0;
            // Q Row 8
            15'b01010001_1000_000: DATA = 1'b1;
            15'b01010001_1000_001: DATA = 1'b1;
            15'b01010001_1000_010: DATA = 1'b0;
            15'b01010001_1000_011: DATA = 1'b0;
            15'b01010001_1000_100: DATA = 1'b0;
            15'b01010001_1000_101: DATA = 1'b1;
            15'b01010001_1000_110: DATA = 1'b1;
            15'b01010001_1000_111: DATA = 1'b0;
            // Q Row 9
            15'b01010001_1001_000: DATA = 1'b1;
            15'b01010001_1001_001: DATA = 1'b1;
            15'b01010001_1001_010: DATA = 1'b0;
            15'b01010001_1001_011: DATA = 1'b1;
            15'b01010001_1001_100: DATA = 1'b0;
            15'b01010001_1001_101: DATA = 1'b1;
            15'b01010001_1001_110: DATA = 1'b1;
            15'b01010001_1001_111: DATA = 1'b0;
            // Q Row 10
            15'b01010001_1010_000: DATA = 1'b1;
            15'b01010001_1010_001: DATA = 1'b1;
            15'b01010001_1010_010: DATA = 1'b0;
            15'b01010001_1010_011: DATA = 1'b0;
            15'b01010001_1010_100: DATA = 1'b1;
            15'b01010001_1010_101: DATA = 1'b1;
            15'b01010001_1010_110: DATA = 1'b1;
            15'b01010001_1010_111: DATA = 1'b0;
            // Q Row 11
            15'b01010001_1011_000: DATA = 1'b0;
            15'b01010001_1011_001: DATA = 1'b1;
            15'b01010001_1011_010: DATA = 1'b1;
            15'b01010001_1011_011: DATA = 1'b1;
            15'b01010001_1011_100: DATA = 1'b1;
            15'b01010001_1011_101: DATA = 1'b1;
            15'b01010001_1011_110: DATA = 1'b0;
            15'b01010001_1011_111: DATA = 1'b0;
            // Q Row 12
            15'b01010001_1100_000: DATA = 1'b0;
            15'b01010001_1100_001: DATA = 1'b0;
            15'b01010001_1100_010: DATA = 1'b1;
            15'b01010001_1100_011: DATA = 1'b1;
            15'b01010001_1100_100: DATA = 1'b1;
            15'b01010001_1100_101: DATA = 1'b0;
            15'b01010001_1100_110: DATA = 1'b1;
            15'b01010001_1100_111: DATA = 1'b0;
            // Q Row 13
            15'b01010001_1101_000: DATA = 1'b0;
            15'b01010001_1101_001: DATA = 1'b0;
            15'b01010001_1101_010: DATA = 1'b0;
            15'b01010001_1101_011: DATA = 1'b0;
            15'b01010001_1101_100: DATA = 1'b0;
            15'b01010001_1101_101: DATA = 1'b0;
            15'b01010001_1101_110: DATA = 1'b0;
            15'b01010001_1101_111: DATA = 1'b0;
            // Q Row 14
            15'b01010001_1110_000: DATA = 1'b0;
            15'b01010001_1110_001: DATA = 1'b0;
            15'b01010001_1110_010: DATA = 1'b0;
            15'b01010001_1110_011: DATA = 1'b0;
            15'b01010001_1110_100: DATA = 1'b0;
            15'b01010001_1110_101: DATA = 1'b0;
            15'b01010001_1110_110: DATA = 1'b0;
            15'b01010001_1110_111: DATA = 1'b0;
            // Q Row 15
            15'b01010001_1111_000: DATA = 1'b0;
            15'b01010001_1111_001: DATA = 1'b0;
            15'b01010001_1111_010: DATA = 1'b0;
            15'b01010001_1111_011: DATA = 1'b0;
            15'b01010001_1111_100: DATA = 1'b0;
            15'b01010001_1111_101: DATA = 1'b0;
            15'b01010001_1111_110: DATA = 1'b0;
            15'b01010001_1111_111: DATA = 1'b0;
            // R Row 0
            15'b01010010_0000_000: DATA = 1'b0;
            15'b01010010_0000_001: DATA = 1'b0;
            15'b01010010_0000_010: DATA = 1'b0;
            15'b01010010_0000_011: DATA = 1'b0;
            15'b01010010_0000_100: DATA = 1'b0;
            15'b01010010_0000_101: DATA = 1'b0;
            15'b01010010_0000_110: DATA = 1'b0;
            15'b01010010_0000_111: DATA = 1'b0;
            // R Row 1
            15'b01010010_0001_000: DATA = 1'b0;
            15'b01010010_0001_001: DATA = 1'b0;
            15'b01010010_0001_010: DATA = 1'b0;
            15'b01010010_0001_011: DATA = 1'b0;
            15'b01010010_0001_100: DATA = 1'b0;
            15'b01010010_0001_101: DATA = 1'b0;
            15'b01010010_0001_110: DATA = 1'b0;
            15'b01010010_0001_111: DATA = 1'b0;
            // R Row 2
            15'b01010010_0010_000: DATA = 1'b0;
            15'b01010010_0010_001: DATA = 1'b0;
            15'b01010010_0010_010: DATA = 1'b0;
            15'b01010010_0010_011: DATA = 1'b0;
            15'b01010010_0010_100: DATA = 1'b0;
            15'b01010010_0010_101: DATA = 1'b0;
            15'b01010010_0010_110: DATA = 1'b0;
            15'b01010010_0010_111: DATA = 1'b0;
            // R Row 3
            15'b01010010_0011_000: DATA = 1'b1;
            15'b01010010_0011_001: DATA = 1'b1;
            15'b01010010_0011_010: DATA = 1'b1;
            15'b01010010_0011_011: DATA = 1'b1;
            15'b01010010_0011_100: DATA = 1'b1;
            15'b01010010_0011_101: DATA = 1'b0;
            15'b01010010_0011_110: DATA = 1'b0;
            15'b01010010_0011_111: DATA = 1'b0;
            // R Row 4
            15'b01010010_0100_000: DATA = 1'b1;
            15'b01010010_0100_001: DATA = 1'b1;
            15'b01010010_0100_010: DATA = 1'b1;
            15'b01010010_0100_011: DATA = 1'b1;
            15'b01010010_0100_100: DATA = 1'b1;
            15'b01010010_0100_101: DATA = 1'b1;
            15'b01010010_0100_110: DATA = 1'b0;
            15'b01010010_0100_111: DATA = 1'b0;
            // R Row 5
            15'b01010010_0101_000: DATA = 1'b1;
            15'b01010010_0101_001: DATA = 1'b1;
            15'b01010010_0101_010: DATA = 1'b0;
            15'b01010010_0101_011: DATA = 1'b0;
            15'b01010010_0101_100: DATA = 1'b0;
            15'b01010010_0101_101: DATA = 1'b1;
            15'b01010010_0101_110: DATA = 1'b1;
            15'b01010010_0101_111: DATA = 1'b0;
            // R Row 6
            15'b01010010_0110_000: DATA = 1'b1;
            15'b01010010_0110_001: DATA = 1'b1;
            15'b01010010_0110_010: DATA = 1'b0;
            15'b01010010_0110_011: DATA = 1'b0;
            15'b01010010_0110_100: DATA = 1'b0;
            15'b01010010_0110_101: DATA = 1'b1;
            15'b01010010_0110_110: DATA = 1'b1;
            15'b01010010_0110_111: DATA = 1'b0;
            // R Row 7
            15'b01010010_0111_000: DATA = 1'b1;
            15'b01010010_0111_001: DATA = 1'b1;
            15'b01010010_0111_010: DATA = 1'b1;
            15'b01010010_0111_011: DATA = 1'b1;
            15'b01010010_0111_100: DATA = 1'b1;
            15'b01010010_0111_101: DATA = 1'b1;
            15'b01010010_0111_110: DATA = 1'b0;
            15'b01010010_0111_111: DATA = 1'b0;
            // R Row 8
            15'b01010010_1000_000: DATA = 1'b1;
            15'b01010010_1000_001: DATA = 1'b1;
            15'b01010010_1000_010: DATA = 1'b1;
            15'b01010010_1000_011: DATA = 1'b1;
            15'b01010010_1000_100: DATA = 1'b1;
            15'b01010010_1000_101: DATA = 1'b0;
            15'b01010010_1000_110: DATA = 1'b0;
            15'b01010010_1000_111: DATA = 1'b0;
            // R Row 9
            15'b01010010_1001_000: DATA = 1'b1;
            15'b01010010_1001_001: DATA = 1'b1;
            15'b01010010_1001_010: DATA = 1'b1;
            15'b01010010_1001_011: DATA = 1'b1;
            15'b01010010_1001_100: DATA = 1'b0;
            15'b01010010_1001_101: DATA = 1'b0;
            15'b01010010_1001_110: DATA = 1'b0;
            15'b01010010_1001_111: DATA = 1'b0;
            // R Row 10
            15'b01010010_1010_000: DATA = 1'b1;
            15'b01010010_1010_001: DATA = 1'b1;
            15'b01010010_1010_010: DATA = 1'b0;
            15'b01010010_1010_011: DATA = 1'b1;
            15'b01010010_1010_100: DATA = 1'b1;
            15'b01010010_1010_101: DATA = 1'b0;
            15'b01010010_1010_110: DATA = 1'b0;
            15'b01010010_1010_111: DATA = 1'b0;
            // R Row 11
            15'b01010010_1011_000: DATA = 1'b1;
            15'b01010010_1011_001: DATA = 1'b1;
            15'b01010010_1011_010: DATA = 1'b0;
            15'b01010010_1011_011: DATA = 1'b0;
            15'b01010010_1011_100: DATA = 1'b1;
            15'b01010010_1011_101: DATA = 1'b1;
            15'b01010010_1011_110: DATA = 1'b0;
            15'b01010010_1011_111: DATA = 1'b0;
            // R Row 12
            15'b01010010_1100_000: DATA = 1'b1;
            15'b01010010_1100_001: DATA = 1'b1;
            15'b01010010_1100_010: DATA = 1'b0;
            15'b01010010_1100_011: DATA = 1'b0;
            15'b01010010_1100_100: DATA = 1'b0;
            15'b01010010_1100_101: DATA = 1'b1;
            15'b01010010_1100_110: DATA = 1'b1;
            15'b01010010_1100_111: DATA = 1'b0;
            // R Row 13
            15'b01010010_1101_000: DATA = 1'b0;
            15'b01010010_1101_001: DATA = 1'b0;
            15'b01010010_1101_010: DATA = 1'b0;
            15'b01010010_1101_011: DATA = 1'b0;
            15'b01010010_1101_100: DATA = 1'b0;
            15'b01010010_1101_101: DATA = 1'b0;
            15'b01010010_1101_110: DATA = 1'b0;
            15'b01010010_1101_111: DATA = 1'b0;
            // R Row 14
            15'b01010010_1110_000: DATA = 1'b0;
            15'b01010010_1110_001: DATA = 1'b0;
            15'b01010010_1110_010: DATA = 1'b0;
            15'b01010010_1110_011: DATA = 1'b0;
            15'b01010010_1110_100: DATA = 1'b0;
            15'b01010010_1110_101: DATA = 1'b0;
            15'b01010010_1110_110: DATA = 1'b0;
            15'b01010010_1110_111: DATA = 1'b0;
            // R Row 15
            15'b01010010_1111_000: DATA = 1'b0;
            15'b01010010_1111_001: DATA = 1'b0;
            15'b01010010_1111_010: DATA = 1'b0;
            15'b01010010_1111_011: DATA = 1'b0;
            15'b01010010_1111_100: DATA = 1'b0;
            15'b01010010_1111_101: DATA = 1'b0;
            15'b01010010_1111_110: DATA = 1'b0;
            15'b01010010_1111_111: DATA = 1'b0;
            // S Row 0
            15'b01010011_0000_000: DATA = 1'b0;
            15'b01010011_0000_001: DATA = 1'b0;
            15'b01010011_0000_010: DATA = 1'b0;
            15'b01010011_0000_011: DATA = 1'b0;
            15'b01010011_0000_100: DATA = 1'b0;
            15'b01010011_0000_101: DATA = 1'b0;
            15'b01010011_0000_110: DATA = 1'b0;
            15'b01010011_0000_111: DATA = 1'b0;
            // S Row 1
            15'b01010011_0001_000: DATA = 1'b0;
            15'b01010011_0001_001: DATA = 1'b0;
            15'b01010011_0001_010: DATA = 1'b0;
            15'b01010011_0001_011: DATA = 1'b0;
            15'b01010011_0001_100: DATA = 1'b0;
            15'b01010011_0001_101: DATA = 1'b0;
            15'b01010011_0001_110: DATA = 1'b0;
            15'b01010011_0001_111: DATA = 1'b0;
            // S Row 2
            15'b01010011_0010_000: DATA = 1'b0;
            15'b01010011_0010_001: DATA = 1'b0;
            15'b01010011_0010_010: DATA = 1'b0;
            15'b01010011_0010_011: DATA = 1'b0;
            15'b01010011_0010_100: DATA = 1'b0;
            15'b01010011_0010_101: DATA = 1'b0;
            15'b01010011_0010_110: DATA = 1'b0;
            15'b01010011_0010_111: DATA = 1'b0;
            // S Row 3
            15'b01010011_0011_000: DATA = 1'b0;
            15'b01010011_0011_001: DATA = 1'b1;
            15'b01010011_0011_010: DATA = 1'b1;
            15'b01010011_0011_011: DATA = 1'b1;
            15'b01010011_0011_100: DATA = 1'b1;
            15'b01010011_0011_101: DATA = 1'b0;
            15'b01010011_0011_110: DATA = 1'b0;
            15'b01010011_0011_111: DATA = 1'b0;
            // S Row 4
            15'b01010011_0100_000: DATA = 1'b1;
            15'b01010011_0100_001: DATA = 1'b1;
            15'b01010011_0100_010: DATA = 1'b0;
            15'b01010011_0100_011: DATA = 1'b0;
            15'b01010011_0100_100: DATA = 1'b1;
            15'b01010011_0100_101: DATA = 1'b1;
            15'b01010011_0100_110: DATA = 1'b0;
            15'b01010011_0100_111: DATA = 1'b0;
            // S Row 5
            15'b01010011_0101_000: DATA = 1'b1;
            15'b01010011_0101_001: DATA = 1'b1;
            15'b01010011_0101_010: DATA = 1'b0;
            15'b01010011_0101_011: DATA = 1'b0;
            15'b01010011_0101_100: DATA = 1'b0;
            15'b01010011_0101_101: DATA = 1'b1;
            15'b01010011_0101_110: DATA = 1'b1;
            15'b01010011_0101_111: DATA = 1'b0;
            // S Row 6
            15'b01010011_0110_000: DATA = 1'b1;
            15'b01010011_0110_001: DATA = 1'b1;
            15'b01010011_0110_010: DATA = 1'b1;
            15'b01010011_0110_011: DATA = 1'b0;
            15'b01010011_0110_100: DATA = 1'b0;
            15'b01010011_0110_101: DATA = 1'b0;
            15'b01010011_0110_110: DATA = 1'b0;
            15'b01010011_0110_111: DATA = 1'b0;
            // S Row 7
            15'b01010011_0111_000: DATA = 1'b0;
            15'b01010011_0111_001: DATA = 1'b1;
            15'b01010011_0111_010: DATA = 1'b1;
            15'b01010011_0111_011: DATA = 1'b1;
            15'b01010011_0111_100: DATA = 1'b1;
            15'b01010011_0111_101: DATA = 1'b1;
            15'b01010011_0111_110: DATA = 1'b0;
            15'b01010011_0111_111: DATA = 1'b0;
            // S Row 8
            15'b01010011_1000_000: DATA = 1'b0;
            15'b01010011_1000_001: DATA = 1'b0;
            15'b01010011_1000_010: DATA = 1'b0;
            15'b01010011_1000_011: DATA = 1'b1;
            15'b01010011_1000_100: DATA = 1'b1;
            15'b01010011_1000_101: DATA = 1'b1;
            15'b01010011_1000_110: DATA = 1'b1;
            15'b01010011_1000_111: DATA = 1'b0;
            // S Row 9
            15'b01010011_1001_000: DATA = 1'b0;
            15'b01010011_1001_001: DATA = 1'b0;
            15'b01010011_1001_010: DATA = 1'b0;
            15'b01010011_1001_011: DATA = 1'b0;
            15'b01010011_1001_100: DATA = 1'b0;
            15'b01010011_1001_101: DATA = 1'b1;
            15'b01010011_1001_110: DATA = 1'b1;
            15'b01010011_1001_111: DATA = 1'b0;
            // S Row 10
            15'b01010011_1010_000: DATA = 1'b1;
            15'b01010011_1010_001: DATA = 1'b1;
            15'b01010011_1010_010: DATA = 1'b0;
            15'b01010011_1010_011: DATA = 1'b0;
            15'b01010011_1010_100: DATA = 1'b0;
            15'b01010011_1010_101: DATA = 1'b1;
            15'b01010011_1010_110: DATA = 1'b1;
            15'b01010011_1010_111: DATA = 1'b0;
            // S Row 11
            15'b01010011_1011_000: DATA = 1'b0;
            15'b01010011_1011_001: DATA = 1'b1;
            15'b01010011_1011_010: DATA = 1'b1;
            15'b01010011_1011_011: DATA = 1'b1;
            15'b01010011_1011_100: DATA = 1'b1;
            15'b01010011_1011_101: DATA = 1'b1;
            15'b01010011_1011_110: DATA = 1'b0;
            15'b01010011_1011_111: DATA = 1'b0;
            // S Row 12
            15'b01010011_1100_000: DATA = 1'b0;
            15'b01010011_1100_001: DATA = 1'b0;
            15'b01010011_1100_010: DATA = 1'b1;
            15'b01010011_1100_011: DATA = 1'b1;
            15'b01010011_1100_100: DATA = 1'b1;
            15'b01010011_1100_101: DATA = 1'b0;
            15'b01010011_1100_110: DATA = 1'b0;
            15'b01010011_1100_111: DATA = 1'b0;
            // S Row 13
            15'b01010011_1101_000: DATA = 1'b0;
            15'b01010011_1101_001: DATA = 1'b0;
            15'b01010011_1101_010: DATA = 1'b0;
            15'b01010011_1101_011: DATA = 1'b0;
            15'b01010011_1101_100: DATA = 1'b0;
            15'b01010011_1101_101: DATA = 1'b0;
            15'b01010011_1101_110: DATA = 1'b0;
            15'b01010011_1101_111: DATA = 1'b0;
            // S Row 14
            15'b01010011_1110_000: DATA = 1'b0;
            15'b01010011_1110_001: DATA = 1'b0;
            15'b01010011_1110_010: DATA = 1'b0;
            15'b01010011_1110_011: DATA = 1'b0;
            15'b01010011_1110_100: DATA = 1'b0;
            15'b01010011_1110_101: DATA = 1'b0;
            15'b01010011_1110_110: DATA = 1'b0;
            15'b01010011_1110_111: DATA = 1'b0;
            // S Row 15
            15'b01010011_1111_000: DATA = 1'b0;
            15'b01010011_1111_001: DATA = 1'b0;
            15'b01010011_1111_010: DATA = 1'b0;
            15'b01010011_1111_011: DATA = 1'b0;
            15'b01010011_1111_100: DATA = 1'b0;
            15'b01010011_1111_101: DATA = 1'b0;
            15'b01010011_1111_110: DATA = 1'b0;
            15'b01010011_1111_111: DATA = 1'b0;
            // T Row 0
            15'b01010100_0000_000: DATA = 1'b0;
            15'b01010100_0000_001: DATA = 1'b0;
            15'b01010100_0000_010: DATA = 1'b0;
            15'b01010100_0000_011: DATA = 1'b0;
            15'b01010100_0000_100: DATA = 1'b0;
            15'b01010100_0000_101: DATA = 1'b0;
            15'b01010100_0000_110: DATA = 1'b0;
            15'b01010100_0000_111: DATA = 1'b0;
            // T Row 1
            15'b01010100_0001_000: DATA = 1'b0;
            15'b01010100_0001_001: DATA = 1'b0;
            15'b01010100_0001_010: DATA = 1'b0;
            15'b01010100_0001_011: DATA = 1'b0;
            15'b01010100_0001_100: DATA = 1'b0;
            15'b01010100_0001_101: DATA = 1'b0;
            15'b01010100_0001_110: DATA = 1'b0;
            15'b01010100_0001_111: DATA = 1'b0;
            // T Row 2
            15'b01010100_0010_000: DATA = 1'b0;
            15'b01010100_0010_001: DATA = 1'b0;
            15'b01010100_0010_010: DATA = 1'b0;
            15'b01010100_0010_011: DATA = 1'b0;
            15'b01010100_0010_100: DATA = 1'b0;
            15'b01010100_0010_101: DATA = 1'b0;
            15'b01010100_0010_110: DATA = 1'b0;
            15'b01010100_0010_111: DATA = 1'b0;
            // T Row 3
            15'b01010100_0011_000: DATA = 1'b1;
            15'b01010100_0011_001: DATA = 1'b1;
            15'b01010100_0011_010: DATA = 1'b1;
            15'b01010100_0011_011: DATA = 1'b1;
            15'b01010100_0011_100: DATA = 1'b1;
            15'b01010100_0011_101: DATA = 1'b1;
            15'b01010100_0011_110: DATA = 1'b1;
            15'b01010100_0011_111: DATA = 1'b0;
            // T Row 4
            15'b01010100_0100_000: DATA = 1'b1;
            15'b01010100_0100_001: DATA = 1'b1;
            15'b01010100_0100_010: DATA = 1'b1;
            15'b01010100_0100_011: DATA = 1'b1;
            15'b01010100_0100_100: DATA = 1'b1;
            15'b01010100_0100_101: DATA = 1'b1;
            15'b01010100_0100_110: DATA = 1'b1;
            15'b01010100_0100_111: DATA = 1'b0;
            // T Row 5
            15'b01010100_0101_000: DATA = 1'b0;
            15'b01010100_0101_001: DATA = 1'b0;
            15'b01010100_0101_010: DATA = 1'b1;
            15'b01010100_0101_011: DATA = 1'b1;
            15'b01010100_0101_100: DATA = 1'b1;
            15'b01010100_0101_101: DATA = 1'b0;
            15'b01010100_0101_110: DATA = 1'b0;
            15'b01010100_0101_111: DATA = 1'b0;
            // T Row 6
            15'b01010100_0110_000: DATA = 1'b0;
            15'b01010100_0110_001: DATA = 1'b0;
            15'b01010100_0110_010: DATA = 1'b1;
            15'b01010100_0110_011: DATA = 1'b1;
            15'b01010100_0110_100: DATA = 1'b1;
            15'b01010100_0110_101: DATA = 1'b0;
            15'b01010100_0110_110: DATA = 1'b0;
            15'b01010100_0110_111: DATA = 1'b0;
            // T Row 7
            15'b01010100_0111_000: DATA = 1'b0;
            15'b01010100_0111_001: DATA = 1'b0;
            15'b01010100_0111_010: DATA = 1'b1;
            15'b01010100_0111_011: DATA = 1'b1;
            15'b01010100_0111_100: DATA = 1'b1;
            15'b01010100_0111_101: DATA = 1'b0;
            15'b01010100_0111_110: DATA = 1'b0;
            15'b01010100_0111_111: DATA = 1'b0;
            // T Row 8
            15'b01010100_1000_000: DATA = 1'b0;
            15'b01010100_1000_001: DATA = 1'b0;
            15'b01010100_1000_010: DATA = 1'b1;
            15'b01010100_1000_011: DATA = 1'b1;
            15'b01010100_1000_100: DATA = 1'b1;
            15'b01010100_1000_101: DATA = 1'b0;
            15'b01010100_1000_110: DATA = 1'b0;
            15'b01010100_1000_111: DATA = 1'b0;
            // T Row 9
            15'b01010100_1001_000: DATA = 1'b0;
            15'b01010100_1001_001: DATA = 1'b0;
            15'b01010100_1001_010: DATA = 1'b1;
            15'b01010100_1001_011: DATA = 1'b1;
            15'b01010100_1001_100: DATA = 1'b1;
            15'b01010100_1001_101: DATA = 1'b0;
            15'b01010100_1001_110: DATA = 1'b0;
            15'b01010100_1001_111: DATA = 1'b0;
            // T Row 10
            15'b01010100_1010_000: DATA = 1'b0;
            15'b01010100_1010_001: DATA = 1'b0;
            15'b01010100_1010_010: DATA = 1'b1;
            15'b01010100_1010_011: DATA = 1'b1;
            15'b01010100_1010_100: DATA = 1'b1;
            15'b01010100_1010_101: DATA = 1'b0;
            15'b01010100_1010_110: DATA = 1'b0;
            15'b01010100_1010_111: DATA = 1'b0;
            // T Row 11
            15'b01010100_1011_000: DATA = 1'b0;
            15'b01010100_1011_001: DATA = 1'b0;
            15'b01010100_1011_010: DATA = 1'b1;
            15'b01010100_1011_011: DATA = 1'b1;
            15'b01010100_1011_100: DATA = 1'b1;
            15'b01010100_1011_101: DATA = 1'b0;
            15'b01010100_1011_110: DATA = 1'b0;
            15'b01010100_1011_111: DATA = 1'b0;
            // T Row 12
            15'b01010100_1100_000: DATA = 1'b0;
            15'b01010100_1100_001: DATA = 1'b0;
            15'b01010100_1100_010: DATA = 1'b1;
            15'b01010100_1100_011: DATA = 1'b1;
            15'b01010100_1100_100: DATA = 1'b1;
            15'b01010100_1100_101: DATA = 1'b0;
            15'b01010100_1100_110: DATA = 1'b0;
            15'b01010100_1100_111: DATA = 1'b0;
            // T Row 13
            15'b01010100_1101_000: DATA = 1'b0;
            15'b01010100_1101_001: DATA = 1'b0;
            15'b01010100_1101_010: DATA = 1'b0;
            15'b01010100_1101_011: DATA = 1'b0;
            15'b01010100_1101_100: DATA = 1'b0;
            15'b01010100_1101_101: DATA = 1'b0;
            15'b01010100_1101_110: DATA = 1'b0;
            15'b01010100_1101_111: DATA = 1'b0;
            // T Row 14
            15'b01010100_1110_000: DATA = 1'b0;
            15'b01010100_1110_001: DATA = 1'b0;
            15'b01010100_1110_010: DATA = 1'b0;
            15'b01010100_1110_011: DATA = 1'b0;
            15'b01010100_1110_100: DATA = 1'b0;
            15'b01010100_1110_101: DATA = 1'b0;
            15'b01010100_1110_110: DATA = 1'b0;
            15'b01010100_1110_111: DATA = 1'b0;
            // T Row 15
            15'b01010100_1111_000: DATA = 1'b0;
            15'b01010100_1111_001: DATA = 1'b0;
            15'b01010100_1111_010: DATA = 1'b0;
            15'b01010100_1111_011: DATA = 1'b0;
            15'b01010100_1111_100: DATA = 1'b0;
            15'b01010100_1111_101: DATA = 1'b0;
            15'b01010100_1111_110: DATA = 1'b0;
            15'b01010100_1111_111: DATA = 1'b0;
            // U Row 0
            15'b01010101_0000_000: DATA = 1'b0;
            15'b01010101_0000_001: DATA = 1'b0;
            15'b01010101_0000_010: DATA = 1'b0;
            15'b01010101_0000_011: DATA = 1'b0;
            15'b01010101_0000_100: DATA = 1'b0;
            15'b01010101_0000_101: DATA = 1'b0;
            15'b01010101_0000_110: DATA = 1'b0;
            15'b01010101_0000_111: DATA = 1'b0;
            // U Row 1
            15'b01010101_0001_000: DATA = 1'b0;
            15'b01010101_0001_001: DATA = 1'b0;
            15'b01010101_0001_010: DATA = 1'b0;
            15'b01010101_0001_011: DATA = 1'b0;
            15'b01010101_0001_100: DATA = 1'b0;
            15'b01010101_0001_101: DATA = 1'b0;
            15'b01010101_0001_110: DATA = 1'b0;
            15'b01010101_0001_111: DATA = 1'b0;
            // U Row 2
            15'b01010101_0010_000: DATA = 1'b0;
            15'b01010101_0010_001: DATA = 1'b0;
            15'b01010101_0010_010: DATA = 1'b0;
            15'b01010101_0010_011: DATA = 1'b0;
            15'b01010101_0010_100: DATA = 1'b0;
            15'b01010101_0010_101: DATA = 1'b0;
            15'b01010101_0010_110: DATA = 1'b0;
            15'b01010101_0010_111: DATA = 1'b0;
            // U Row 3
            15'b01010101_0011_000: DATA = 1'b1;
            15'b01010101_0011_001: DATA = 1'b1;
            15'b01010101_0011_010: DATA = 1'b0;
            15'b01010101_0011_011: DATA = 1'b0;
            15'b01010101_0011_100: DATA = 1'b0;
            15'b01010101_0011_101: DATA = 1'b0;
            15'b01010101_0011_110: DATA = 1'b1;
            15'b01010101_0011_111: DATA = 1'b0;
            // U Row 4
            15'b01010101_0100_000: DATA = 1'b1;
            15'b01010101_0100_001: DATA = 1'b1;
            15'b01010101_0100_010: DATA = 1'b0;
            15'b01010101_0100_011: DATA = 1'b0;
            15'b01010101_0100_100: DATA = 1'b0;
            15'b01010101_0100_101: DATA = 1'b0;
            15'b01010101_0100_110: DATA = 1'b1;
            15'b01010101_0100_111: DATA = 1'b0;
            // U Row 5
            15'b01010101_0101_000: DATA = 1'b1;
            15'b01010101_0101_001: DATA = 1'b1;
            15'b01010101_0101_010: DATA = 1'b0;
            15'b01010101_0101_011: DATA = 1'b0;
            15'b01010101_0101_100: DATA = 1'b0;
            15'b01010101_0101_101: DATA = 1'b0;
            15'b01010101_0101_110: DATA = 1'b1;
            15'b01010101_0101_111: DATA = 1'b0;
            // U Row 6
            15'b01010101_0110_000: DATA = 1'b1;
            15'b01010101_0110_001: DATA = 1'b1;
            15'b01010101_0110_010: DATA = 1'b0;
            15'b01010101_0110_011: DATA = 1'b0;
            15'b01010101_0110_100: DATA = 1'b0;
            15'b01010101_0110_101: DATA = 1'b0;
            15'b01010101_0110_110: DATA = 1'b1;
            15'b01010101_0110_111: DATA = 1'b0;
            // U Row 7
            15'b01010101_0111_000: DATA = 1'b1;
            15'b01010101_0111_001: DATA = 1'b1;
            15'b01010101_0111_010: DATA = 1'b0;
            15'b01010101_0111_011: DATA = 1'b0;
            15'b01010101_0111_100: DATA = 1'b0;
            15'b01010101_0111_101: DATA = 1'b0;
            15'b01010101_0111_110: DATA = 1'b1;
            15'b01010101_0111_111: DATA = 1'b0;
            // U Row 8
            15'b01010101_1000_000: DATA = 1'b1;
            15'b01010101_1000_001: DATA = 1'b1;
            15'b01010101_1000_010: DATA = 1'b0;
            15'b01010101_1000_011: DATA = 1'b0;
            15'b01010101_1000_100: DATA = 1'b0;
            15'b01010101_1000_101: DATA = 1'b0;
            15'b01010101_1000_110: DATA = 1'b1;
            15'b01010101_1000_111: DATA = 1'b0;
            // U Row 9
            15'b01010101_1001_000: DATA = 1'b1;
            15'b01010101_1001_001: DATA = 1'b1;
            15'b01010101_1001_010: DATA = 1'b0;
            15'b01010101_1001_011: DATA = 1'b0;
            15'b01010101_1001_100: DATA = 1'b0;
            15'b01010101_1001_101: DATA = 1'b0;
            15'b01010101_1001_110: DATA = 1'b1;
            15'b01010101_1001_111: DATA = 1'b0;
            // U Row 10
            15'b01010101_1010_000: DATA = 1'b0;
            15'b01010101_1010_001: DATA = 1'b1;
            15'b01010101_1010_010: DATA = 1'b1;
            15'b01010101_1010_011: DATA = 1'b0;
            15'b01010101_1010_100: DATA = 1'b0;
            15'b01010101_1010_101: DATA = 1'b0;
            15'b01010101_1010_110: DATA = 1'b1;
            15'b01010101_1010_111: DATA = 1'b0;
            // U Row 11
            15'b01010101_1011_000: DATA = 1'b0;
            15'b01010101_1011_001: DATA = 1'b1;
            15'b01010101_1011_010: DATA = 1'b1;
            15'b01010101_1011_011: DATA = 1'b1;
            15'b01010101_1011_100: DATA = 1'b0;
            15'b01010101_1011_101: DATA = 1'b1;
            15'b01010101_1011_110: DATA = 1'b1;
            15'b01010101_1011_111: DATA = 1'b0;
            // U Row 12
            15'b01010101_1100_000: DATA = 1'b0;
            15'b01010101_1100_001: DATA = 1'b0;
            15'b01010101_1100_010: DATA = 1'b1;
            15'b01010101_1100_011: DATA = 1'b1;
            15'b01010101_1100_100: DATA = 1'b1;
            15'b01010101_1100_101: DATA = 1'b1;
            15'b01010101_1100_110: DATA = 1'b0;
            15'b01010101_1100_111: DATA = 1'b0;
            // U Row 13
            15'b01010101_1101_000: DATA = 1'b0;
            15'b01010101_1101_001: DATA = 1'b0;
            15'b01010101_1101_010: DATA = 1'b0;
            15'b01010101_1101_011: DATA = 1'b0;
            15'b01010101_1101_100: DATA = 1'b0;
            15'b01010101_1101_101: DATA = 1'b0;
            15'b01010101_1101_110: DATA = 1'b0;
            15'b01010101_1101_111: DATA = 1'b0;
            // U Row 14
            15'b01010101_1110_000: DATA = 1'b0;
            15'b01010101_1110_001: DATA = 1'b0;
            15'b01010101_1110_010: DATA = 1'b0;
            15'b01010101_1110_011: DATA = 1'b0;
            15'b01010101_1110_100: DATA = 1'b0;
            15'b01010101_1110_101: DATA = 1'b0;
            15'b01010101_1110_110: DATA = 1'b0;
            15'b01010101_1110_111: DATA = 1'b0;
            // U Row 15
            15'b01010101_1111_000: DATA = 1'b0;
            15'b01010101_1111_001: DATA = 1'b0;
            15'b01010101_1111_010: DATA = 1'b0;
            15'b01010101_1111_011: DATA = 1'b0;
            15'b01010101_1111_100: DATA = 1'b0;
            15'b01010101_1111_101: DATA = 1'b0;
            15'b01010101_1111_110: DATA = 1'b0;
            15'b01010101_1111_111: DATA = 1'b0;
            // V Row 0
            15'b01010110_0000_000: DATA = 1'b0;
            15'b01010110_0000_001: DATA = 1'b0;
            15'b01010110_0000_010: DATA = 1'b0;
            15'b01010110_0000_011: DATA = 1'b0;
            15'b01010110_0000_100: DATA = 1'b0;
            15'b01010110_0000_101: DATA = 1'b0;
            15'b01010110_0000_110: DATA = 1'b0;
            15'b01010110_0000_111: DATA = 1'b0;
            // V Row 1
            15'b01010110_0001_000: DATA = 1'b0;
            15'b01010110_0001_001: DATA = 1'b0;
            15'b01010110_0001_010: DATA = 1'b0;
            15'b01010110_0001_011: DATA = 1'b0;
            15'b01010110_0001_100: DATA = 1'b0;
            15'b01010110_0001_101: DATA = 1'b0;
            15'b01010110_0001_110: DATA = 1'b0;
            15'b01010110_0001_111: DATA = 1'b0;
            // V Row 2
            15'b01010110_0010_000: DATA = 1'b0;
            15'b01010110_0010_001: DATA = 1'b0;
            15'b01010110_0010_010: DATA = 1'b0;
            15'b01010110_0010_011: DATA = 1'b0;
            15'b01010110_0010_100: DATA = 1'b0;
            15'b01010110_0010_101: DATA = 1'b0;
            15'b01010110_0010_110: DATA = 1'b0;
            15'b01010110_0010_111: DATA = 1'b0;
            // V Row 3
            15'b01010110_0011_000: DATA = 1'b1;
            15'b01010110_0011_001: DATA = 1'b1;
            15'b01010110_0011_010: DATA = 1'b0;
            15'b01010110_0011_011: DATA = 1'b0;
            15'b01010110_0011_100: DATA = 1'b0;
            15'b01010110_0011_101: DATA = 1'b0;
            15'b01010110_0011_110: DATA = 1'b1;
            15'b01010110_0011_111: DATA = 1'b0;
            // V Row 4
            15'b01010110_0100_000: DATA = 1'b1;
            15'b01010110_0100_001: DATA = 1'b1;
            15'b01010110_0100_010: DATA = 1'b0;
            15'b01010110_0100_011: DATA = 1'b0;
            15'b01010110_0100_100: DATA = 1'b0;
            15'b01010110_0100_101: DATA = 1'b0;
            15'b01010110_0100_110: DATA = 1'b1;
            15'b01010110_0100_111: DATA = 1'b0;
            // V Row 5
            15'b01010110_0101_000: DATA = 1'b1;
            15'b01010110_0101_001: DATA = 1'b1;
            15'b01010110_0101_010: DATA = 1'b0;
            15'b01010110_0101_011: DATA = 1'b0;
            15'b01010110_0101_100: DATA = 1'b0;
            15'b01010110_0101_101: DATA = 1'b0;
            15'b01010110_0101_110: DATA = 1'b1;
            15'b01010110_0101_111: DATA = 1'b0;
            // V Row 6
            15'b01010110_0110_000: DATA = 1'b0;
            15'b01010110_0110_001: DATA = 1'b1;
            15'b01010110_0110_010: DATA = 1'b1;
            15'b01010110_0110_011: DATA = 1'b0;
            15'b01010110_0110_100: DATA = 1'b0;
            15'b01010110_0110_101: DATA = 1'b0;
            15'b01010110_0110_110: DATA = 1'b1;
            15'b01010110_0110_111: DATA = 1'b0;
            // V Row 7
            15'b01010110_0111_000: DATA = 1'b0;
            15'b01010110_0111_001: DATA = 1'b1;
            15'b01010110_0111_010: DATA = 1'b1;
            15'b01010110_0111_011: DATA = 1'b0;
            15'b01010110_0111_100: DATA = 1'b0;
            15'b01010110_0111_101: DATA = 1'b1;
            15'b01010110_0111_110: DATA = 1'b1;
            15'b01010110_0111_111: DATA = 1'b0;
            // V Row 8
            15'b01010110_1000_000: DATA = 1'b0;
            15'b01010110_1000_001: DATA = 1'b0;
            15'b01010110_1000_010: DATA = 1'b1;
            15'b01010110_1000_011: DATA = 1'b0;
            15'b01010110_1000_100: DATA = 1'b0;
            15'b01010110_1000_101: DATA = 1'b1;
            15'b01010110_1000_110: DATA = 1'b0;
            15'b01010110_1000_111: DATA = 1'b0;
            // V Row 9
            15'b01010110_1001_000: DATA = 1'b0;
            15'b01010110_1001_001: DATA = 1'b0;
            15'b01010110_1001_010: DATA = 1'b1;
            15'b01010110_1001_011: DATA = 1'b1;
            15'b01010110_1001_100: DATA = 1'b0;
            15'b01010110_1001_101: DATA = 1'b1;
            15'b01010110_1001_110: DATA = 1'b0;
            15'b01010110_1001_111: DATA = 1'b0;
            // V Row 10
            15'b01010110_1010_000: DATA = 1'b0;
            15'b01010110_1010_001: DATA = 1'b0;
            15'b01010110_1010_010: DATA = 1'b1;
            15'b01010110_1010_011: DATA = 1'b1;
            15'b01010110_1010_100: DATA = 1'b0;
            15'b01010110_1010_101: DATA = 1'b1;
            15'b01010110_1010_110: DATA = 1'b0;
            15'b01010110_1010_111: DATA = 1'b0;
            // V Row 11
            15'b01010110_1011_000: DATA = 1'b0;
            15'b01010110_1011_001: DATA = 1'b0;
            15'b01010110_1011_010: DATA = 1'b0;
            15'b01010110_1011_011: DATA = 1'b1;
            15'b01010110_1011_100: DATA = 1'b1;
            15'b01010110_1011_101: DATA = 1'b0;
            15'b01010110_1011_110: DATA = 1'b0;
            15'b01010110_1011_111: DATA = 1'b0;
            // V Row 12
            15'b01010110_1100_000: DATA = 1'b0;
            15'b01010110_1100_001: DATA = 1'b0;
            15'b01010110_1100_010: DATA = 1'b0;
            15'b01010110_1100_011: DATA = 1'b1;
            15'b01010110_1100_100: DATA = 1'b1;
            15'b01010110_1100_101: DATA = 1'b0;
            15'b01010110_1100_110: DATA = 1'b0;
            15'b01010110_1100_111: DATA = 1'b0;
            // V Row 13
            15'b01010110_1101_000: DATA = 1'b0;
            15'b01010110_1101_001: DATA = 1'b0;
            15'b01010110_1101_010: DATA = 1'b0;
            15'b01010110_1101_011: DATA = 1'b0;
            15'b01010110_1101_100: DATA = 1'b0;
            15'b01010110_1101_101: DATA = 1'b0;
            15'b01010110_1101_110: DATA = 1'b0;
            15'b01010110_1101_111: DATA = 1'b0;
            // V Row 14
            15'b01010110_1110_000: DATA = 1'b0;
            15'b01010110_1110_001: DATA = 1'b0;
            15'b01010110_1110_010: DATA = 1'b0;
            15'b01010110_1110_011: DATA = 1'b0;
            15'b01010110_1110_100: DATA = 1'b0;
            15'b01010110_1110_101: DATA = 1'b0;
            15'b01010110_1110_110: DATA = 1'b0;
            15'b01010110_1110_111: DATA = 1'b0;
            // V Row 15
            15'b01010110_1111_000: DATA = 1'b0;
            15'b01010110_1111_001: DATA = 1'b0;
            15'b01010110_1111_010: DATA = 1'b0;
            15'b01010110_1111_011: DATA = 1'b0;
            15'b01010110_1111_100: DATA = 1'b0;
            15'b01010110_1111_101: DATA = 1'b0;
            15'b01010110_1111_110: DATA = 1'b0;
            15'b01010110_1111_111: DATA = 1'b0;
            // W Row 0
            15'b01010111_0000_000: DATA = 1'b0;
            15'b01010111_0000_001: DATA = 1'b0;
            15'b01010111_0000_010: DATA = 1'b0;
            15'b01010111_0000_011: DATA = 1'b0;
            15'b01010111_0000_100: DATA = 1'b0;
            15'b01010111_0000_101: DATA = 1'b0;
            15'b01010111_0000_110: DATA = 1'b0;
            15'b01010111_0000_111: DATA = 1'b0;
            // W Row 1
            15'b01010111_0001_000: DATA = 1'b0;
            15'b01010111_0001_001: DATA = 1'b0;
            15'b01010111_0001_010: DATA = 1'b0;
            15'b01010111_0001_011: DATA = 1'b0;
            15'b01010111_0001_100: DATA = 1'b0;
            15'b01010111_0001_101: DATA = 1'b0;
            15'b01010111_0001_110: DATA = 1'b0;
            15'b01010111_0001_111: DATA = 1'b0;
            // W Row 2
            15'b01010111_0010_000: DATA = 1'b0;
            15'b01010111_0010_001: DATA = 1'b0;
            15'b01010111_0010_010: DATA = 1'b0;
            15'b01010111_0010_011: DATA = 1'b0;
            15'b01010111_0010_100: DATA = 1'b0;
            15'b01010111_0010_101: DATA = 1'b0;
            15'b01010111_0010_110: DATA = 1'b0;
            15'b01010111_0010_111: DATA = 1'b0;
            // W Row 3
            15'b01010111_0011_000: DATA = 1'b1;
            15'b01010111_0011_001: DATA = 1'b1;
            15'b01010111_0011_010: DATA = 1'b0;
            15'b01010111_0011_011: DATA = 1'b0;
            15'b01010111_0011_100: DATA = 1'b0;
            15'b01010111_0011_101: DATA = 1'b0;
            15'b01010111_0011_110: DATA = 1'b1;
            15'b01010111_0011_111: DATA = 1'b0;
            // W Row 4
            15'b01010111_0100_000: DATA = 1'b1;
            15'b01010111_0100_001: DATA = 1'b1;
            15'b01010111_0100_010: DATA = 1'b0;
            15'b01010111_0100_011: DATA = 1'b0;
            15'b01010111_0100_100: DATA = 1'b0;
            15'b01010111_0100_101: DATA = 1'b0;
            15'b01010111_0100_110: DATA = 1'b1;
            15'b01010111_0100_111: DATA = 1'b0;
            // W Row 5
            15'b01010111_0101_000: DATA = 1'b1;
            15'b01010111_0101_001: DATA = 1'b1;
            15'b01010111_0101_010: DATA = 1'b0;
            15'b01010111_0101_011: DATA = 1'b0;
            15'b01010111_0101_100: DATA = 1'b0;
            15'b01010111_0101_101: DATA = 1'b0;
            15'b01010111_0101_110: DATA = 1'b1;
            15'b01010111_0101_111: DATA = 1'b0;
            // W Row 6
            15'b01010111_0110_000: DATA = 1'b1;
            15'b01010111_0110_001: DATA = 1'b1;
            15'b01010111_0110_010: DATA = 1'b0;
            15'b01010111_0110_011: DATA = 1'b0;
            15'b01010111_0110_100: DATA = 1'b0;
            15'b01010111_0110_101: DATA = 1'b0;
            15'b01010111_0110_110: DATA = 1'b1;
            15'b01010111_0110_111: DATA = 1'b0;
            // W Row 7
            15'b01010111_0111_000: DATA = 1'b1;
            15'b01010111_0111_001: DATA = 1'b1;
            15'b01010111_0111_010: DATA = 1'b0;
            15'b01010111_0111_011: DATA = 1'b0;
            15'b01010111_0111_100: DATA = 1'b1;
            15'b01010111_0111_101: DATA = 1'b0;
            15'b01010111_0111_110: DATA = 1'b1;
            15'b01010111_0111_111: DATA = 1'b0;
            // W Row 8
            15'b01010111_1000_000: DATA = 1'b1;
            15'b01010111_1000_001: DATA = 1'b1;
            15'b01010111_1000_010: DATA = 1'b0;
            15'b01010111_1000_011: DATA = 1'b0;
            15'b01010111_1000_100: DATA = 1'b1;
            15'b01010111_1000_101: DATA = 1'b0;
            15'b01010111_1000_110: DATA = 1'b1;
            15'b01010111_1000_111: DATA = 1'b0;
            // W Row 9
            15'b01010111_1001_000: DATA = 1'b1;
            15'b01010111_1001_001: DATA = 1'b1;
            15'b01010111_1001_010: DATA = 1'b0;
            15'b01010111_1001_011: DATA = 1'b0;
            15'b01010111_1001_100: DATA = 1'b1;
            15'b01010111_1001_101: DATA = 1'b0;
            15'b01010111_1001_110: DATA = 1'b1;
            15'b01010111_1001_111: DATA = 1'b0;
            // W Row 10
            15'b01010111_1010_000: DATA = 1'b1;
            15'b01010111_1010_001: DATA = 1'b1;
            15'b01010111_1010_010: DATA = 1'b0;
            15'b01010111_1010_011: DATA = 1'b1;
            15'b01010111_1010_100: DATA = 1'b1;
            15'b01010111_1010_101: DATA = 1'b0;
            15'b01010111_1010_110: DATA = 1'b1;
            15'b01010111_1010_111: DATA = 1'b0;
            // W Row 11
            15'b01010111_1011_000: DATA = 1'b0;
            15'b01010111_1011_001: DATA = 1'b1;
            15'b01010111_1011_010: DATA = 1'b1;
            15'b01010111_1011_011: DATA = 1'b1;
            15'b01010111_1011_100: DATA = 1'b1;
            15'b01010111_1011_101: DATA = 1'b1;
            15'b01010111_1011_110: DATA = 1'b1;
            15'b01010111_1011_111: DATA = 1'b0;
            // W Row 12
            15'b01010111_1100_000: DATA = 1'b0;
            15'b01010111_1100_001: DATA = 1'b0;
            15'b01010111_1100_010: DATA = 1'b1;
            15'b01010111_1100_011: DATA = 1'b1;
            15'b01010111_1100_100: DATA = 1'b1;
            15'b01010111_1100_101: DATA = 1'b1;
            15'b01010111_1100_110: DATA = 1'b0;
            15'b01010111_1100_111: DATA = 1'b0;
            // W Row 13
            15'b01010111_1101_000: DATA = 1'b0;
            15'b01010111_1101_001: DATA = 1'b0;
            15'b01010111_1101_010: DATA = 1'b0;
            15'b01010111_1101_011: DATA = 1'b0;
            15'b01010111_1101_100: DATA = 1'b0;
            15'b01010111_1101_101: DATA = 1'b0;
            15'b01010111_1101_110: DATA = 1'b0;
            15'b01010111_1101_111: DATA = 1'b0;
            // W Row 14
            15'b01010111_1110_000: DATA = 1'b0;
            15'b01010111_1110_001: DATA = 1'b0;
            15'b01010111_1110_010: DATA = 1'b0;
            15'b01010111_1110_011: DATA = 1'b0;
            15'b01010111_1110_100: DATA = 1'b0;
            15'b01010111_1110_101: DATA = 1'b0;
            15'b01010111_1110_110: DATA = 1'b0;
            15'b01010111_1110_111: DATA = 1'b0;
            // W Row 15
            15'b01010111_1111_000: DATA = 1'b0;
            15'b01010111_1111_001: DATA = 1'b0;
            15'b01010111_1111_010: DATA = 1'b0;
            15'b01010111_1111_011: DATA = 1'b0;
            15'b01010111_1111_100: DATA = 1'b0;
            15'b01010111_1111_101: DATA = 1'b0;
            15'b01010111_1111_110: DATA = 1'b0;
            15'b01010111_1111_111: DATA = 1'b0;
            // X Row 0
            15'b01011000_0000_000: DATA = 1'b0;
            15'b01011000_0000_001: DATA = 1'b0;
            15'b01011000_0000_010: DATA = 1'b0;
            15'b01011000_0000_011: DATA = 1'b0;
            15'b01011000_0000_100: DATA = 1'b0;
            15'b01011000_0000_101: DATA = 1'b0;
            15'b01011000_0000_110: DATA = 1'b0;
            15'b01011000_0000_111: DATA = 1'b0;
            // X Row 1
            15'b01011000_0001_000: DATA = 1'b0;
            15'b01011000_0001_001: DATA = 1'b0;
            15'b01011000_0001_010: DATA = 1'b0;
            15'b01011000_0001_011: DATA = 1'b0;
            15'b01011000_0001_100: DATA = 1'b0;
            15'b01011000_0001_101: DATA = 1'b0;
            15'b01011000_0001_110: DATA = 1'b0;
            15'b01011000_0001_111: DATA = 1'b0;
            // X Row 2
            15'b01011000_0010_000: DATA = 1'b0;
            15'b01011000_0010_001: DATA = 1'b0;
            15'b01011000_0010_010: DATA = 1'b0;
            15'b01011000_0010_011: DATA = 1'b0;
            15'b01011000_0010_100: DATA = 1'b0;
            15'b01011000_0010_101: DATA = 1'b0;
            15'b01011000_0010_110: DATA = 1'b0;
            15'b01011000_0010_111: DATA = 1'b0;
            // X Row 3
            15'b01011000_0011_000: DATA = 1'b1;
            15'b01011000_0011_001: DATA = 1'b1;
            15'b01011000_0011_010: DATA = 1'b0;
            15'b01011000_0011_011: DATA = 1'b0;
            15'b01011000_0011_100: DATA = 1'b0;
            15'b01011000_0011_101: DATA = 1'b1;
            15'b01011000_0011_110: DATA = 1'b1;
            15'b01011000_0011_111: DATA = 1'b0;
            // X Row 4
            15'b01011000_0100_000: DATA = 1'b0;
            15'b01011000_0100_001: DATA = 1'b1;
            15'b01011000_0100_010: DATA = 1'b0;
            15'b01011000_0100_011: DATA = 1'b0;
            15'b01011000_0100_100: DATA = 1'b0;
            15'b01011000_0100_101: DATA = 1'b1;
            15'b01011000_0100_110: DATA = 1'b0;
            15'b01011000_0100_111: DATA = 1'b0;
            // X Row 5
            15'b01011000_0101_000: DATA = 1'b0;
            15'b01011000_0101_001: DATA = 1'b1;
            15'b01011000_0101_010: DATA = 1'b1;
            15'b01011000_0101_011: DATA = 1'b0;
            15'b01011000_0101_100: DATA = 1'b1;
            15'b01011000_0101_101: DATA = 1'b1;
            15'b01011000_0101_110: DATA = 1'b0;
            15'b01011000_0101_111: DATA = 1'b0;
            // X Row 6
            15'b01011000_0110_000: DATA = 1'b0;
            15'b01011000_0110_001: DATA = 1'b1;
            15'b01011000_0110_010: DATA = 1'b1;
            15'b01011000_0110_011: DATA = 1'b1;
            15'b01011000_0110_100: DATA = 1'b1;
            15'b01011000_0110_101: DATA = 1'b1;
            15'b01011000_0110_110: DATA = 1'b0;
            15'b01011000_0110_111: DATA = 1'b0;
            // X Row 7
            15'b01011000_0111_000: DATA = 1'b0;
            15'b01011000_0111_001: DATA = 1'b0;
            15'b01011000_0111_010: DATA = 1'b1;
            15'b01011000_0111_011: DATA = 1'b1;
            15'b01011000_0111_100: DATA = 1'b1;
            15'b01011000_0111_101: DATA = 1'b0;
            15'b01011000_0111_110: DATA = 1'b0;
            15'b01011000_0111_111: DATA = 1'b0;
            // X Row 8
            15'b01011000_1000_000: DATA = 1'b0;
            15'b01011000_1000_001: DATA = 1'b0;
            15'b01011000_1000_010: DATA = 1'b1;
            15'b01011000_1000_011: DATA = 1'b1;
            15'b01011000_1000_100: DATA = 1'b1;
            15'b01011000_1000_101: DATA = 1'b0;
            15'b01011000_1000_110: DATA = 1'b0;
            15'b01011000_1000_111: DATA = 1'b0;
            // X Row 9
            15'b01011000_1001_000: DATA = 1'b0;
            15'b01011000_1001_001: DATA = 1'b1;
            15'b01011000_1001_010: DATA = 1'b1;
            15'b01011000_1001_011: DATA = 1'b1;
            15'b01011000_1001_100: DATA = 1'b1;
            15'b01011000_1001_101: DATA = 1'b1;
            15'b01011000_1001_110: DATA = 1'b0;
            15'b01011000_1001_111: DATA = 1'b0;
            // X Row 10
            15'b01011000_1010_000: DATA = 1'b0;
            15'b01011000_1010_001: DATA = 1'b1;
            15'b01011000_1010_010: DATA = 1'b1;
            15'b01011000_1010_011: DATA = 1'b0;
            15'b01011000_1010_100: DATA = 1'b1;
            15'b01011000_1010_101: DATA = 1'b1;
            15'b01011000_1010_110: DATA = 1'b0;
            15'b01011000_1010_111: DATA = 1'b0;
            // X Row 11
            15'b01011000_1011_000: DATA = 1'b0;
            15'b01011000_1011_001: DATA = 1'b1;
            15'b01011000_1011_010: DATA = 1'b0;
            15'b01011000_1011_011: DATA = 1'b0;
            15'b01011000_1011_100: DATA = 1'b0;
            15'b01011000_1011_101: DATA = 1'b1;
            15'b01011000_1011_110: DATA = 1'b0;
            15'b01011000_1011_111: DATA = 1'b0;
            // X Row 12
            15'b01011000_1100_000: DATA = 1'b1;
            15'b01011000_1100_001: DATA = 1'b1;
            15'b01011000_1100_010: DATA = 1'b0;
            15'b01011000_1100_011: DATA = 1'b0;
            15'b01011000_1100_100: DATA = 1'b0;
            15'b01011000_1100_101: DATA = 1'b1;
            15'b01011000_1100_110: DATA = 1'b1;
            15'b01011000_1100_111: DATA = 1'b0;
            // X Row 13
            15'b01011000_1101_000: DATA = 1'b0;
            15'b01011000_1101_001: DATA = 1'b0;
            15'b01011000_1101_010: DATA = 1'b0;
            15'b01011000_1101_011: DATA = 1'b0;
            15'b01011000_1101_100: DATA = 1'b0;
            15'b01011000_1101_101: DATA = 1'b0;
            15'b01011000_1101_110: DATA = 1'b0;
            15'b01011000_1101_111: DATA = 1'b0;
            // X Row 14
            15'b01011000_1110_000: DATA = 1'b0;
            15'b01011000_1110_001: DATA = 1'b0;
            15'b01011000_1110_010: DATA = 1'b0;
            15'b01011000_1110_011: DATA = 1'b0;
            15'b01011000_1110_100: DATA = 1'b0;
            15'b01011000_1110_101: DATA = 1'b0;
            15'b01011000_1110_110: DATA = 1'b0;
            15'b01011000_1110_111: DATA = 1'b0;
            // X Row 15
            15'b01011000_1111_000: DATA = 1'b0;
            15'b01011000_1111_001: DATA = 1'b0;
            15'b01011000_1111_010: DATA = 1'b0;
            15'b01011000_1111_011: DATA = 1'b0;
            15'b01011000_1111_100: DATA = 1'b0;
            15'b01011000_1111_101: DATA = 1'b0;
            15'b01011000_1111_110: DATA = 1'b0;
            15'b01011000_1111_111: DATA = 1'b0;
            // Y Row 0
            15'b01011001_0000_000: DATA = 1'b0;
            15'b01011001_0000_001: DATA = 1'b0;
            15'b01011001_0000_010: DATA = 1'b0;
            15'b01011001_0000_011: DATA = 1'b0;
            15'b01011001_0000_100: DATA = 1'b0;
            15'b01011001_0000_101: DATA = 1'b0;
            15'b01011001_0000_110: DATA = 1'b0;
            15'b01011001_0000_111: DATA = 1'b0;
            // Y Row 1
            15'b01011001_0001_000: DATA = 1'b0;
            15'b01011001_0001_001: DATA = 1'b0;
            15'b01011001_0001_010: DATA = 1'b0;
            15'b01011001_0001_011: DATA = 1'b0;
            15'b01011001_0001_100: DATA = 1'b0;
            15'b01011001_0001_101: DATA = 1'b0;
            15'b01011001_0001_110: DATA = 1'b0;
            15'b01011001_0001_111: DATA = 1'b0;
            // Y Row 2
            15'b01011001_0010_000: DATA = 1'b0;
            15'b01011001_0010_001: DATA = 1'b0;
            15'b01011001_0010_010: DATA = 1'b0;
            15'b01011001_0010_011: DATA = 1'b0;
            15'b01011001_0010_100: DATA = 1'b0;
            15'b01011001_0010_101: DATA = 1'b0;
            15'b01011001_0010_110: DATA = 1'b0;
            15'b01011001_0010_111: DATA = 1'b0;
            // Y Row 3
            15'b01011001_0011_000: DATA = 1'b1;
            15'b01011001_0011_001: DATA = 1'b1;
            15'b01011001_0011_010: DATA = 1'b0;
            15'b01011001_0011_011: DATA = 1'b0;
            15'b01011001_0011_100: DATA = 1'b0;
            15'b01011001_0011_101: DATA = 1'b1;
            15'b01011001_0011_110: DATA = 1'b1;
            15'b01011001_0011_111: DATA = 1'b0;
            // Y Row 4
            15'b01011001_0100_000: DATA = 1'b1;
            15'b01011001_0100_001: DATA = 1'b1;
            15'b01011001_0100_010: DATA = 1'b0;
            15'b01011001_0100_011: DATA = 1'b0;
            15'b01011001_0100_100: DATA = 1'b0;
            15'b01011001_0100_101: DATA = 1'b1;
            15'b01011001_0100_110: DATA = 1'b1;
            15'b01011001_0100_111: DATA = 1'b0;
            // Y Row 5
            15'b01011001_0101_000: DATA = 1'b1;
            15'b01011001_0101_001: DATA = 1'b1;
            15'b01011001_0101_010: DATA = 1'b0;
            15'b01011001_0101_011: DATA = 1'b0;
            15'b01011001_0101_100: DATA = 1'b0;
            15'b01011001_0101_101: DATA = 1'b1;
            15'b01011001_0101_110: DATA = 1'b1;
            15'b01011001_0101_111: DATA = 1'b0;
            // Y Row 6
            15'b01011001_0110_000: DATA = 1'b1;
            15'b01011001_0110_001: DATA = 1'b1;
            15'b01011001_0110_010: DATA = 1'b0;
            15'b01011001_0110_011: DATA = 1'b0;
            15'b01011001_0110_100: DATA = 1'b0;
            15'b01011001_0110_101: DATA = 1'b1;
            15'b01011001_0110_110: DATA = 1'b1;
            15'b01011001_0110_111: DATA = 1'b0;
            // Y Row 7
            15'b01011001_0111_000: DATA = 1'b0;
            15'b01011001_0111_001: DATA = 1'b1;
            15'b01011001_0111_010: DATA = 1'b1;
            15'b01011001_0111_011: DATA = 1'b1;
            15'b01011001_0111_100: DATA = 1'b1;
            15'b01011001_0111_101: DATA = 1'b1;
            15'b01011001_0111_110: DATA = 1'b0;
            15'b01011001_0111_111: DATA = 1'b0;
            // Y Row 8
            15'b01011001_1000_000: DATA = 1'b0;
            15'b01011001_1000_001: DATA = 1'b0;
            15'b01011001_1000_010: DATA = 1'b1;
            15'b01011001_1000_011: DATA = 1'b1;
            15'b01011001_1000_100: DATA = 1'b1;
            15'b01011001_1000_101: DATA = 1'b0;
            15'b01011001_1000_110: DATA = 1'b0;
            15'b01011001_1000_111: DATA = 1'b0;
            // Y Row 9
            15'b01011001_1001_000: DATA = 1'b0;
            15'b01011001_1001_001: DATA = 1'b0;
            15'b01011001_1001_010: DATA = 1'b1;
            15'b01011001_1001_011: DATA = 1'b1;
            15'b01011001_1001_100: DATA = 1'b1;
            15'b01011001_1001_101: DATA = 1'b0;
            15'b01011001_1001_110: DATA = 1'b0;
            15'b01011001_1001_111: DATA = 1'b0;
            // Y Row 10
            15'b01011001_1010_000: DATA = 1'b0;
            15'b01011001_1010_001: DATA = 1'b0;
            15'b01011001_1010_010: DATA = 1'b1;
            15'b01011001_1010_011: DATA = 1'b1;
            15'b01011001_1010_100: DATA = 1'b1;
            15'b01011001_1010_101: DATA = 1'b0;
            15'b01011001_1010_110: DATA = 1'b0;
            15'b01011001_1010_111: DATA = 1'b0;
            // Y Row 11
            15'b01011001_1011_000: DATA = 1'b0;
            15'b01011001_1011_001: DATA = 1'b0;
            15'b01011001_1011_010: DATA = 1'b1;
            15'b01011001_1011_011: DATA = 1'b1;
            15'b01011001_1011_100: DATA = 1'b1;
            15'b01011001_1011_101: DATA = 1'b0;
            15'b01011001_1011_110: DATA = 1'b0;
            15'b01011001_1011_111: DATA = 1'b0;
            // Y Row 12
            15'b01011001_1100_000: DATA = 1'b0;
            15'b01011001_1100_001: DATA = 1'b0;
            15'b01011001_1100_010: DATA = 1'b1;
            15'b01011001_1100_011: DATA = 1'b1;
            15'b01011001_1100_100: DATA = 1'b1;
            15'b01011001_1100_101: DATA = 1'b0;
            15'b01011001_1100_110: DATA = 1'b0;
            15'b01011001_1100_111: DATA = 1'b0;
            // Y Row 13
            15'b01011001_1101_000: DATA = 1'b0;
            15'b01011001_1101_001: DATA = 1'b0;
            15'b01011001_1101_010: DATA = 1'b0;
            15'b01011001_1101_011: DATA = 1'b0;
            15'b01011001_1101_100: DATA = 1'b0;
            15'b01011001_1101_101: DATA = 1'b0;
            15'b01011001_1101_110: DATA = 1'b0;
            15'b01011001_1101_111: DATA = 1'b0;
            // Y Row 14
            15'b01011001_1110_000: DATA = 1'b0;
            15'b01011001_1110_001: DATA = 1'b0;
            15'b01011001_1110_010: DATA = 1'b0;
            15'b01011001_1110_011: DATA = 1'b0;
            15'b01011001_1110_100: DATA = 1'b0;
            15'b01011001_1110_101: DATA = 1'b0;
            15'b01011001_1110_110: DATA = 1'b0;
            15'b01011001_1110_111: DATA = 1'b0;
            // Y Row 15
            15'b01011001_1111_000: DATA = 1'b0;
            15'b01011001_1111_001: DATA = 1'b0;
            15'b01011001_1111_010: DATA = 1'b0;
            15'b01011001_1111_011: DATA = 1'b0;
            15'b01011001_1111_100: DATA = 1'b0;
            15'b01011001_1111_101: DATA = 1'b0;
            15'b01011001_1111_110: DATA = 1'b0;
            15'b01011001_1111_111: DATA = 1'b0;
            // Z Row 0
            15'b01011010_0000_000: DATA = 1'b0;
            15'b01011010_0000_001: DATA = 1'b0;
            15'b01011010_0000_010: DATA = 1'b0;
            15'b01011010_0000_011: DATA = 1'b0;
            15'b01011010_0000_100: DATA = 1'b0;
            15'b01011010_0000_101: DATA = 1'b0;
            15'b01011010_0000_110: DATA = 1'b0;
            15'b01011010_0000_111: DATA = 1'b0;
            // Z Row 1
            15'b01011010_0001_000: DATA = 1'b0;
            15'b01011010_0001_001: DATA = 1'b0;
            15'b01011010_0001_010: DATA = 1'b0;
            15'b01011010_0001_011: DATA = 1'b0;
            15'b01011010_0001_100: DATA = 1'b0;
            15'b01011010_0001_101: DATA = 1'b0;
            15'b01011010_0001_110: DATA = 1'b0;
            15'b01011010_0001_111: DATA = 1'b0;
            // Z Row 2
            15'b01011010_0010_000: DATA = 1'b0;
            15'b01011010_0010_001: DATA = 1'b0;
            15'b01011010_0010_010: DATA = 1'b0;
            15'b01011010_0010_011: DATA = 1'b0;
            15'b01011010_0010_100: DATA = 1'b0;
            15'b01011010_0010_101: DATA = 1'b0;
            15'b01011010_0010_110: DATA = 1'b0;
            15'b01011010_0010_111: DATA = 1'b0;
            // Z Row 3
            15'b01011010_0011_000: DATA = 1'b1;
            15'b01011010_0011_001: DATA = 1'b1;
            15'b01011010_0011_010: DATA = 1'b1;
            15'b01011010_0011_011: DATA = 1'b1;
            15'b01011010_0011_100: DATA = 1'b1;
            15'b01011010_0011_101: DATA = 1'b1;
            15'b01011010_0011_110: DATA = 1'b1;
            15'b01011010_0011_111: DATA = 1'b0;
            // Z Row 4
            15'b01011010_0100_000: DATA = 1'b1;
            15'b01011010_0100_001: DATA = 1'b1;
            15'b01011010_0100_010: DATA = 1'b1;
            15'b01011010_0100_011: DATA = 1'b1;
            15'b01011010_0100_100: DATA = 1'b1;
            15'b01011010_0100_101: DATA = 1'b1;
            15'b01011010_0100_110: DATA = 1'b1;
            15'b01011010_0100_111: DATA = 1'b0;
            // Z Row 5
            15'b01011010_0101_000: DATA = 1'b0;
            15'b01011010_0101_001: DATA = 1'b0;
            15'b01011010_0101_010: DATA = 1'b0;
            15'b01011010_0101_011: DATA = 1'b0;
            15'b01011010_0101_100: DATA = 1'b0;
            15'b01011010_0101_101: DATA = 1'b1;
            15'b01011010_0101_110: DATA = 1'b1;
            15'b01011010_0101_111: DATA = 1'b0;
            // Z Row 6
            15'b01011010_0110_000: DATA = 1'b0;
            15'b01011010_0110_001: DATA = 1'b0;
            15'b01011010_0110_010: DATA = 1'b0;
            15'b01011010_0110_011: DATA = 1'b0;
            15'b01011010_0110_100: DATA = 1'b1;
            15'b01011010_0110_101: DATA = 1'b1;
            15'b01011010_0110_110: DATA = 1'b0;
            15'b01011010_0110_111: DATA = 1'b0;
            // Z Row 7
            15'b01011010_0111_000: DATA = 1'b0;
            15'b01011010_0111_001: DATA = 1'b0;
            15'b01011010_0111_010: DATA = 1'b0;
            15'b01011010_0111_011: DATA = 1'b1;
            15'b01011010_0111_100: DATA = 1'b1;
            15'b01011010_0111_101: DATA = 1'b0;
            15'b01011010_0111_110: DATA = 1'b0;
            15'b01011010_0111_111: DATA = 1'b0;
            // Z Row 8
            15'b01011010_1000_000: DATA = 1'b0;
            15'b01011010_1000_001: DATA = 1'b0;
            15'b01011010_1000_010: DATA = 1'b1;
            15'b01011010_1000_011: DATA = 1'b1;
            15'b01011010_1000_100: DATA = 1'b0;
            15'b01011010_1000_101: DATA = 1'b0;
            15'b01011010_1000_110: DATA = 1'b0;
            15'b01011010_1000_111: DATA = 1'b0;
            // Z Row 9
            15'b01011010_1001_000: DATA = 1'b0;
            15'b01011010_1001_001: DATA = 1'b1;
            15'b01011010_1001_010: DATA = 1'b1;
            15'b01011010_1001_011: DATA = 1'b0;
            15'b01011010_1001_100: DATA = 1'b0;
            15'b01011010_1001_101: DATA = 1'b0;
            15'b01011010_1001_110: DATA = 1'b0;
            15'b01011010_1001_111: DATA = 1'b0;
            // Z Row 10
            15'b01011010_1010_000: DATA = 1'b1;
            15'b01011010_1010_001: DATA = 1'b1;
            15'b01011010_1010_010: DATA = 1'b0;
            15'b01011010_1010_011: DATA = 1'b0;
            15'b01011010_1010_100: DATA = 1'b0;
            15'b01011010_1010_101: DATA = 1'b0;
            15'b01011010_1010_110: DATA = 1'b0;
            15'b01011010_1010_111: DATA = 1'b0;
            // Z Row 11
            15'b01011010_1011_000: DATA = 1'b1;
            15'b01011010_1011_001: DATA = 1'b1;
            15'b01011010_1011_010: DATA = 1'b1;
            15'b01011010_1011_011: DATA = 1'b1;
            15'b01011010_1011_100: DATA = 1'b1;
            15'b01011010_1011_101: DATA = 1'b1;
            15'b01011010_1011_110: DATA = 1'b1;
            15'b01011010_1011_111: DATA = 1'b0;
            // Z Row 12
            15'b01011010_1100_000: DATA = 1'b1;
            15'b01011010_1100_001: DATA = 1'b1;
            15'b01011010_1100_010: DATA = 1'b1;
            15'b01011010_1100_011: DATA = 1'b1;
            15'b01011010_1100_100: DATA = 1'b1;
            15'b01011010_1100_101: DATA = 1'b1;
            15'b01011010_1100_110: DATA = 1'b1;
            15'b01011010_1100_111: DATA = 1'b0;
            // Z Row 13
            15'b01011010_1101_000: DATA = 1'b0;
            15'b01011010_1101_001: DATA = 1'b0;
            15'b01011010_1101_010: DATA = 1'b0;
            15'b01011010_1101_011: DATA = 1'b0;
            15'b01011010_1101_100: DATA = 1'b0;
            15'b01011010_1101_101: DATA = 1'b0;
            15'b01011010_1101_110: DATA = 1'b0;
            15'b01011010_1101_111: DATA = 1'b0;
            // Z Row 14
            15'b01011010_1110_000: DATA = 1'b0;
            15'b01011010_1110_001: DATA = 1'b0;
            15'b01011010_1110_010: DATA = 1'b0;
            15'b01011010_1110_011: DATA = 1'b0;
            15'b01011010_1110_100: DATA = 1'b0;
            15'b01011010_1110_101: DATA = 1'b0;
            15'b01011010_1110_110: DATA = 1'b0;
            15'b01011010_1110_111: DATA = 1'b0;
            // Z Row 15
            15'b01011010_1111_000: DATA = 1'b0;
            15'b01011010_1111_001: DATA = 1'b0;
            15'b01011010_1111_010: DATA = 1'b0;
            15'b01011010_1111_011: DATA = 1'b0;
            15'b01011010_1111_100: DATA = 1'b0;
            15'b01011010_1111_101: DATA = 1'b0;
            15'b01011010_1111_110: DATA = 1'b0;
            15'b01011010_1111_111: DATA = 1'b0;
            
            
            // PICTURES
            // SINE+ ROW 0 COL 0 Row 0
            15'b10000000_0000_000: DATA = 1'b0;
            15'b10000000_0000_001: DATA = 1'b0;
            15'b10000000_0000_010: DATA = 1'b0;
            15'b10000000_0000_011: DATA = 1'b0;
            15'b10000000_0000_100: DATA = 1'b0;
            15'b10000000_0000_101: DATA = 1'b0;
            15'b10000000_0000_110: DATA = 1'b0;
            15'b10000000_0000_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 0 Row 1
            15'b10000000_0001_000: DATA = 1'b0;
            15'b10000000_0001_001: DATA = 1'b0;
            15'b10000000_0001_010: DATA = 1'b0;
            15'b10000000_0001_011: DATA = 1'b0;
            15'b10000000_0001_100: DATA = 1'b0;
            15'b10000000_0001_101: DATA = 1'b0;
            15'b10000000_0001_110: DATA = 1'b0;
            15'b10000000_0001_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 0 Row 2
            15'b10000000_0010_000: DATA = 1'b0;
            15'b10000000_0010_001: DATA = 1'b0;
            15'b10000000_0010_010: DATA = 1'b0;
            15'b10000000_0010_011: DATA = 1'b0;
            15'b10000000_0010_100: DATA = 1'b0;
            15'b10000000_0010_101: DATA = 1'b0;
            15'b10000000_0010_110: DATA = 1'b0;
            15'b10000000_0010_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 0 Row 3
            15'b10000000_0011_000: DATA = 1'b0;
            15'b10000000_0011_001: DATA = 1'b0;
            15'b10000000_0011_010: DATA = 1'b0;
            15'b10000000_0011_011: DATA = 1'b0;
            15'b10000000_0011_100: DATA = 1'b0;
            15'b10000000_0011_101: DATA = 1'b0;
            15'b10000000_0011_110: DATA = 1'b0;
            15'b10000000_0011_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 0 Row 4
            15'b10000000_0100_000: DATA = 1'b0;
            15'b10000000_0100_001: DATA = 1'b0;
            15'b10000000_0100_010: DATA = 1'b0;
            15'b10000000_0100_011: DATA = 1'b0;
            15'b10000000_0100_100: DATA = 1'b0;
            15'b10000000_0100_101: DATA = 1'b0;
            15'b10000000_0100_110: DATA = 1'b0;
            15'b10000000_0100_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 0 Row 5
            15'b10000000_0101_000: DATA = 1'b0;
            15'b10000000_0101_001: DATA = 1'b0;
            15'b10000000_0101_010: DATA = 1'b0;
            15'b10000000_0101_011: DATA = 1'b0;
            15'b10000000_0101_100: DATA = 1'b0;
            15'b10000000_0101_101: DATA = 1'b0;
            15'b10000000_0101_110: DATA = 1'b0;
            15'b10000000_0101_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 0 Row 6
            15'b10000000_0110_000: DATA = 1'b0;
            15'b10000000_0110_001: DATA = 1'b0;
            15'b10000000_0110_010: DATA = 1'b0;
            15'b10000000_0110_011: DATA = 1'b0;
            15'b10000000_0110_100: DATA = 1'b0;
            15'b10000000_0110_101: DATA = 1'b0;
            15'b10000000_0110_110: DATA = 1'b0;
            15'b10000000_0110_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 0 Row 7
            15'b10000000_0111_000: DATA = 1'b0;
            15'b10000000_0111_001: DATA = 1'b0;
            15'b10000000_0111_010: DATA = 1'b0;
            15'b10000000_0111_011: DATA = 1'b0;
            15'b10000000_0111_100: DATA = 1'b0;
            15'b10000000_0111_101: DATA = 1'b0;
            15'b10000000_0111_110: DATA = 1'b0;
            15'b10000000_0111_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 0 Row 8
            15'b10000000_1000_000: DATA = 1'b0;
            15'b10000000_1000_001: DATA = 1'b0;
            15'b10000000_1000_010: DATA = 1'b0;
            15'b10000000_1000_011: DATA = 1'b0;
            15'b10000000_1000_100: DATA = 1'b0;
            15'b10000000_1000_101: DATA = 1'b0;
            15'b10000000_1000_110: DATA = 1'b0;
            15'b10000000_1000_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 0 Row 9
            15'b10000000_1001_000: DATA = 1'b0;
            15'b10000000_1001_001: DATA = 1'b0;
            15'b10000000_1001_010: DATA = 1'b0;
            15'b10000000_1001_011: DATA = 1'b0;
            15'b10000000_1001_100: DATA = 1'b0;
            15'b10000000_1001_101: DATA = 1'b0;
            15'b10000000_1001_110: DATA = 1'b0;
            15'b10000000_1001_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 0 Row 10
            15'b10000000_1010_000: DATA = 1'b0;
            15'b10000000_1010_001: DATA = 1'b0;
            15'b10000000_1010_010: DATA = 1'b0;
            15'b10000000_1010_011: DATA = 1'b0;
            15'b10000000_1010_100: DATA = 1'b0;
            15'b10000000_1010_101: DATA = 1'b0;
            15'b10000000_1010_110: DATA = 1'b0;
            15'b10000000_1010_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 0 Row 11
            15'b10000000_1011_000: DATA = 1'b0;
            15'b10000000_1011_001: DATA = 1'b0;
            15'b10000000_1011_010: DATA = 1'b0;
            15'b10000000_1011_011: DATA = 1'b0;
            15'b10000000_1011_100: DATA = 1'b0;
            15'b10000000_1011_101: DATA = 1'b0;
            15'b10000000_1011_110: DATA = 1'b0;
            15'b10000000_1011_111: DATA = 1'b1;
            // SINE+ ROW 0 COL 0 Row 12
            15'b10000000_1100_000: DATA = 1'b0;
            15'b10000000_1100_001: DATA = 1'b0;
            15'b10000000_1100_010: DATA = 1'b0;
            15'b10000000_1100_011: DATA = 1'b0;
            15'b10000000_1100_100: DATA = 1'b0;
            15'b10000000_1100_101: DATA = 1'b0;
            15'b10000000_1100_110: DATA = 1'b0;
            15'b10000000_1100_111: DATA = 1'b1;
            // SINE+ ROW 0 COL 0 Row 13
            15'b10000000_1101_000: DATA = 1'b0;
            15'b10000000_1101_001: DATA = 1'b0;
            15'b10000000_1101_010: DATA = 1'b0;
            15'b10000000_1101_011: DATA = 1'b0;
            15'b10000000_1101_100: DATA = 1'b0;
            15'b10000000_1101_101: DATA = 1'b0;
            15'b10000000_1101_110: DATA = 1'b1;
            15'b10000000_1101_111: DATA = 1'b1;
            // SINE+ ROW 0 COL 0 Row 14
            15'b10000000_1110_000: DATA = 1'b0;
            15'b10000000_1110_001: DATA = 1'b0;
            15'b10000000_1110_010: DATA = 1'b0;
            15'b10000000_1110_011: DATA = 1'b0;
            15'b10000000_1110_100: DATA = 1'b0;
            15'b10000000_1110_101: DATA = 1'b0;
            15'b10000000_1110_110: DATA = 1'b1;
            15'b10000000_1110_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 0 Row 15
            15'b10000000_1111_000: DATA = 1'b0;
            15'b10000000_1111_001: DATA = 1'b0;
            15'b10000000_1111_010: DATA = 1'b0;
            15'b10000000_1111_011: DATA = 1'b0;
            15'b10000000_1111_100: DATA = 1'b0;
            15'b10000000_1111_101: DATA = 1'b1;
            15'b10000000_1111_110: DATA = 1'b1;
            15'b10000000_1111_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 1 Row 0
            15'b10000001_0000_000: DATA = 1'b0;
            15'b10000001_0000_001: DATA = 1'b0;
            15'b10000001_0000_010: DATA = 1'b0;
            15'b10000001_0000_011: DATA = 1'b0;
            15'b10000001_0000_100: DATA = 1'b0;
            15'b10000001_0000_101: DATA = 1'b0;
            15'b10000001_0000_110: DATA = 1'b0;
            15'b10000001_0000_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 1 Row 1
            15'b10000001_0001_000: DATA = 1'b0;
            15'b10000001_0001_001: DATA = 1'b0;
            15'b10000001_0001_010: DATA = 1'b0;
            15'b10000001_0001_011: DATA = 1'b0;
            15'b10000001_0001_100: DATA = 1'b0;
            15'b10000001_0001_101: DATA = 1'b0;
            15'b10000001_0001_110: DATA = 1'b0;
            15'b10000001_0001_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 1 Row 2
            15'b10000001_0010_000: DATA = 1'b0;
            15'b10000001_0010_001: DATA = 1'b0;
            15'b10000001_0010_010: DATA = 1'b0;
            15'b10000001_0010_011: DATA = 1'b0;
            15'b10000001_0010_100: DATA = 1'b0;
            15'b10000001_0010_101: DATA = 1'b0;
            15'b10000001_0010_110: DATA = 1'b1;
            15'b10000001_0010_111: DATA = 1'b1;
            // SINE+ ROW 0 COL 1 Row 3
            15'b10000001_0011_000: DATA = 1'b0;
            15'b10000001_0011_001: DATA = 1'b0;
            15'b10000001_0011_010: DATA = 1'b0;
            15'b10000001_0011_011: DATA = 1'b0;
            15'b10000001_0011_100: DATA = 1'b0;
            15'b10000001_0011_101: DATA = 1'b1;
            15'b10000001_0011_110: DATA = 1'b1;
            15'b10000001_0011_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 1 Row 4
            15'b10000001_0100_000: DATA = 1'b0;
            15'b10000001_0100_001: DATA = 1'b0;
            15'b10000001_0100_010: DATA = 1'b0;
            15'b10000001_0100_011: DATA = 1'b0;
            15'b10000001_0100_100: DATA = 1'b1;
            15'b10000001_0100_101: DATA = 1'b1;
            15'b10000001_0100_110: DATA = 1'b0;
            15'b10000001_0100_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 1 Row 5
            15'b10000001_0101_000: DATA = 1'b0;
            15'b10000001_0101_001: DATA = 1'b0;
            15'b10000001_0101_010: DATA = 1'b0;
            15'b10000001_0101_011: DATA = 1'b1;
            15'b10000001_0101_100: DATA = 1'b1;
            15'b10000001_0101_101: DATA = 1'b0;
            15'b10000001_0101_110: DATA = 1'b0;
            15'b10000001_0101_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 1 Row 6
            15'b10000001_0110_000: DATA = 1'b0;
            15'b10000001_0110_001: DATA = 1'b0;
            15'b10000001_0110_010: DATA = 1'b1;
            15'b10000001_0110_011: DATA = 1'b1;
            15'b10000001_0110_100: DATA = 1'b0;
            15'b10000001_0110_101: DATA = 1'b0;
            15'b10000001_0110_110: DATA = 1'b0;
            15'b10000001_0110_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 1 Row 7
            15'b10000001_0111_000: DATA = 1'b0;
            15'b10000001_0111_001: DATA = 1'b1;
            15'b10000001_0111_010: DATA = 1'b1;
            15'b10000001_0111_011: DATA = 1'b0;
            15'b10000001_0111_100: DATA = 1'b0;
            15'b10000001_0111_101: DATA = 1'b0;
            15'b10000001_0111_110: DATA = 1'b0;
            15'b10000001_0111_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 1 Row 8
            15'b10000001_1000_000: DATA = 1'b0;
            15'b10000001_1000_001: DATA = 1'b1;
            15'b10000001_1000_010: DATA = 1'b0;
            15'b10000001_1000_011: DATA = 1'b0;
            15'b10000001_1000_100: DATA = 1'b0;
            15'b10000001_1000_101: DATA = 1'b0;
            15'b10000001_1000_110: DATA = 1'b0;
            15'b10000001_1000_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 1 Row 9
            15'b10000001_1001_000: DATA = 1'b1;
            15'b10000001_1001_001: DATA = 1'b1;
            15'b10000001_1001_010: DATA = 1'b0;
            15'b10000001_1001_011: DATA = 1'b0;
            15'b10000001_1001_100: DATA = 1'b0;
            15'b10000001_1001_101: DATA = 1'b0;
            15'b10000001_1001_110: DATA = 1'b0;
            15'b10000001_1001_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 1 Row 10
            15'b10000001_1010_000: DATA = 1'b1;
            15'b10000001_1010_001: DATA = 1'b0;
            15'b10000001_1010_010: DATA = 1'b0;
            15'b10000001_1010_011: DATA = 1'b0;
            15'b10000001_1010_100: DATA = 1'b0;
            15'b10000001_1010_101: DATA = 1'b0;
            15'b10000001_1010_110: DATA = 1'b0;
            15'b10000001_1010_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 1 Row 11
            15'b10000001_1011_000: DATA = 1'b1;
            15'b10000001_1011_001: DATA = 1'b0;
            15'b10000001_1011_010: DATA = 1'b0;
            15'b10000001_1011_011: DATA = 1'b0;
            15'b10000001_1011_100: DATA = 1'b0;
            15'b10000001_1011_101: DATA = 1'b0;
            15'b10000001_1011_110: DATA = 1'b0;
            15'b10000001_1011_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 1 Row 12
            15'b10000001_1100_000: DATA = 1'b0;
            15'b10000001_1100_001: DATA = 1'b0;
            15'b10000001_1100_010: DATA = 1'b0;
            15'b10000001_1100_011: DATA = 1'b0;
            15'b10000001_1100_100: DATA = 1'b0;
            15'b10000001_1100_101: DATA = 1'b0;
            15'b10000001_1100_110: DATA = 1'b0;
            15'b10000001_1100_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 1 Row 13
            15'b10000001_1101_000: DATA = 1'b0;
            15'b10000001_1101_001: DATA = 1'b0;
            15'b10000001_1101_010: DATA = 1'b0;
            15'b10000001_1101_011: DATA = 1'b0;
            15'b10000001_1101_100: DATA = 1'b0;
            15'b10000001_1101_101: DATA = 1'b0;
            15'b10000001_1101_110: DATA = 1'b0;
            15'b10000001_1101_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 1 Row 14
            15'b10000001_1110_000: DATA = 1'b0;
            15'b10000001_1110_001: DATA = 1'b0;
            15'b10000001_1110_010: DATA = 1'b0;
            15'b10000001_1110_011: DATA = 1'b0;
            15'b10000001_1110_100: DATA = 1'b0;
            15'b10000001_1110_101: DATA = 1'b0;
            15'b10000001_1110_110: DATA = 1'b0;
            15'b10000001_1110_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 1 Row 15
            15'b10000001_1111_000: DATA = 1'b0;
            15'b10000001_1111_001: DATA = 1'b0;
            15'b10000001_1111_010: DATA = 1'b0;
            15'b10000001_1111_011: DATA = 1'b0;
            15'b10000001_1111_100: DATA = 1'b0;
            15'b10000001_1111_101: DATA = 1'b0;
            15'b10000001_1111_110: DATA = 1'b0;
            15'b10000001_1111_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 2 Row 0
            15'b10000010_0000_000: DATA = 1'b0;
            15'b10000010_0000_001: DATA = 1'b0;
            15'b10000010_0000_010: DATA = 1'b1;
            15'b10000010_0000_011: DATA = 1'b1;
            15'b10000010_0000_100: DATA = 1'b1;
            15'b10000010_0000_101: DATA = 1'b1;
            15'b10000010_0000_110: DATA = 1'b0;
            15'b10000010_0000_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 2 Row 1
            15'b10000010_0001_000: DATA = 1'b1;
            15'b10000010_0001_001: DATA = 1'b1;
            15'b10000010_0001_010: DATA = 1'b1;
            15'b10000010_0001_011: DATA = 1'b0;
            15'b10000010_0001_100: DATA = 1'b0;
            15'b10000010_0001_101: DATA = 1'b1;
            15'b10000010_0001_110: DATA = 1'b1;
            15'b10000010_0001_111: DATA = 1'b1;
            // SINE+ ROW 0 COL 2 Row 2
            15'b10000010_0010_000: DATA = 1'b1;
            15'b10000010_0010_001: DATA = 1'b0;
            15'b10000010_0010_010: DATA = 1'b0;
            15'b10000010_0010_011: DATA = 1'b0;
            15'b10000010_0010_100: DATA = 1'b0;
            15'b10000010_0010_101: DATA = 1'b0;
            15'b10000010_0010_110: DATA = 1'b0;
            15'b10000010_0010_111: DATA = 1'b1;
            // SINE+ ROW 0 COL 2 Row 3
            15'b10000010_0011_000: DATA = 1'b0;
            15'b10000010_0011_001: DATA = 1'b0;
            15'b10000010_0011_010: DATA = 1'b0;
            15'b10000010_0011_011: DATA = 1'b0;
            15'b10000010_0011_100: DATA = 1'b0;
            15'b10000010_0011_101: DATA = 1'b0;
            15'b10000010_0011_110: DATA = 1'b0;
            15'b10000010_0011_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 2 Row 4
            15'b10000010_0100_000: DATA = 1'b0;
            15'b10000010_0100_001: DATA = 1'b0;
            15'b10000010_0100_010: DATA = 1'b0;
            15'b10000010_0100_011: DATA = 1'b0;
            15'b10000010_0100_100: DATA = 1'b0;
            15'b10000010_0100_101: DATA = 1'b0;
            15'b10000010_0100_110: DATA = 1'b0;
            15'b10000010_0100_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 2 Row 5
            15'b10000010_0101_000: DATA = 1'b0;
            15'b10000010_0101_001: DATA = 1'b0;
            15'b10000010_0101_010: DATA = 1'b0;
            15'b10000010_0101_011: DATA = 1'b0;
            15'b10000010_0101_100: DATA = 1'b0;
            15'b10000010_0101_101: DATA = 1'b0;
            15'b10000010_0101_110: DATA = 1'b0;
            15'b10000010_0101_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 2 Row 6
            15'b10000010_0110_000: DATA = 1'b0;
            15'b10000010_0110_001: DATA = 1'b0;
            15'b10000010_0110_010: DATA = 1'b0;
            15'b10000010_0110_011: DATA = 1'b0;
            15'b10000010_0110_100: DATA = 1'b0;
            15'b10000010_0110_101: DATA = 1'b0;
            15'b10000010_0110_110: DATA = 1'b0;
            15'b10000010_0110_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 2 Row 7
            15'b10000010_0111_000: DATA = 1'b0;
            15'b10000010_0111_001: DATA = 1'b0;
            15'b10000010_0111_010: DATA = 1'b0;
            15'b10000010_0111_011: DATA = 1'b0;
            15'b10000010_0111_100: DATA = 1'b0;
            15'b10000010_0111_101: DATA = 1'b0;
            15'b10000010_0111_110: DATA = 1'b0;
            15'b10000010_0111_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 2 Row 8
            15'b10000010_1000_000: DATA = 1'b0;
            15'b10000010_1000_001: DATA = 1'b0;
            15'b10000010_1000_010: DATA = 1'b0;
            15'b10000010_1000_011: DATA = 1'b0;
            15'b10000010_1000_100: DATA = 1'b0;
            15'b10000010_1000_101: DATA = 1'b0;
            15'b10000010_1000_110: DATA = 1'b0;
            15'b10000010_1000_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 2 Row 9
            15'b10000010_1001_000: DATA = 1'b0;
            15'b10000010_1001_001: DATA = 1'b0;
            15'b10000010_1001_010: DATA = 1'b0;
            15'b10000010_1001_011: DATA = 1'b0;
            15'b10000010_1001_100: DATA = 1'b0;
            15'b10000010_1001_101: DATA = 1'b0;
            15'b10000010_1001_110: DATA = 1'b0;
            15'b10000010_1001_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 2 Row 10
            15'b10000010_1010_000: DATA = 1'b0;
            15'b10000010_1010_001: DATA = 1'b0;
            15'b10000010_1010_010: DATA = 1'b0;
            15'b10000010_1010_011: DATA = 1'b0;
            15'b10000010_1010_100: DATA = 1'b0;
            15'b10000010_1010_101: DATA = 1'b0;
            15'b10000010_1010_110: DATA = 1'b0;
            15'b10000010_1010_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 2 Row 11
            15'b10000010_1011_000: DATA = 1'b0;
            15'b10000010_1011_001: DATA = 1'b0;
            15'b10000010_1011_010: DATA = 1'b0;
            15'b10000010_1011_011: DATA = 1'b0;
            15'b10000010_1011_100: DATA = 1'b0;
            15'b10000010_1011_101: DATA = 1'b0;
            15'b10000010_1011_110: DATA = 1'b0;
            15'b10000010_1011_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 2 Row 12
            15'b10000010_1100_000: DATA = 1'b0;
            15'b10000010_1100_001: DATA = 1'b0;
            15'b10000010_1100_010: DATA = 1'b0;
            15'b10000010_1100_011: DATA = 1'b0;
            15'b10000010_1100_100: DATA = 1'b0;
            15'b10000010_1100_101: DATA = 1'b0;
            15'b10000010_1100_110: DATA = 1'b0;
            15'b10000010_1100_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 2 Row 13
            15'b10000010_1101_000: DATA = 1'b0;
            15'b10000010_1101_001: DATA = 1'b0;
            15'b10000010_1101_010: DATA = 1'b0;
            15'b10000010_1101_011: DATA = 1'b0;
            15'b10000010_1101_100: DATA = 1'b0;
            15'b10000010_1101_101: DATA = 1'b0;
            15'b10000010_1101_110: DATA = 1'b0;
            15'b10000010_1101_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 2 Row 14
            15'b10000010_1110_000: DATA = 1'b0;
            15'b10000010_1110_001: DATA = 1'b0;
            15'b10000010_1110_010: DATA = 1'b0;
            15'b10000010_1110_011: DATA = 1'b0;
            15'b10000010_1110_100: DATA = 1'b0;
            15'b10000010_1110_101: DATA = 1'b0;
            15'b10000010_1110_110: DATA = 1'b0;
            15'b10000010_1110_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 2 Row 15
            15'b10000010_1111_000: DATA = 1'b0;
            15'b10000010_1111_001: DATA = 1'b0;
            15'b10000010_1111_010: DATA = 1'b0;
            15'b10000010_1111_011: DATA = 1'b0;
            15'b10000010_1111_100: DATA = 1'b0;
            15'b10000010_1111_101: DATA = 1'b0;
            15'b10000010_1111_110: DATA = 1'b0;
            15'b10000010_1111_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 3 Row 0
            15'b10000011_0000_000: DATA = 1'b0;
            15'b10000011_0000_001: DATA = 1'b0;
            15'b10000011_0000_010: DATA = 1'b0;
            15'b10000011_0000_011: DATA = 1'b0;
            15'b10000011_0000_100: DATA = 1'b0;
            15'b10000011_0000_101: DATA = 1'b0;
            15'b10000011_0000_110: DATA = 1'b0;
            15'b10000011_0000_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 3 Row 1
            15'b10000011_0001_000: DATA = 1'b0;
            15'b10000011_0001_001: DATA = 1'b0;
            15'b10000011_0001_010: DATA = 1'b0;
            15'b10000011_0001_011: DATA = 1'b0;
            15'b10000011_0001_100: DATA = 1'b0;
            15'b10000011_0001_101: DATA = 1'b0;
            15'b10000011_0001_110: DATA = 1'b0;
            15'b10000011_0001_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 3 Row 2
            15'b10000011_0010_000: DATA = 1'b1;
            15'b10000011_0010_001: DATA = 1'b1;
            15'b10000011_0010_010: DATA = 1'b0;
            15'b10000011_0010_011: DATA = 1'b0;
            15'b10000011_0010_100: DATA = 1'b0;
            15'b10000011_0010_101: DATA = 1'b0;
            15'b10000011_0010_110: DATA = 1'b0;
            15'b10000011_0010_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 3 Row 3
            15'b10000011_0011_000: DATA = 1'b0;
            15'b10000011_0011_001: DATA = 1'b1;
            15'b10000011_0011_010: DATA = 1'b1;
            15'b10000011_0011_011: DATA = 1'b0;
            15'b10000011_0011_100: DATA = 1'b0;
            15'b10000011_0011_101: DATA = 1'b0;
            15'b10000011_0011_110: DATA = 1'b0;
            15'b10000011_0011_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 3 Row 4
            15'b10000011_0100_000: DATA = 1'b0;
            15'b10000011_0100_001: DATA = 1'b0;
            15'b10000011_0100_010: DATA = 1'b1;
            15'b10000011_0100_011: DATA = 1'b1;
            15'b10000011_0100_100: DATA = 1'b0;
            15'b10000011_0100_101: DATA = 1'b0;
            15'b10000011_0100_110: DATA = 1'b0;
            15'b10000011_0100_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 3 Row 5
            15'b10000011_0101_000: DATA = 1'b0;
            15'b10000011_0101_001: DATA = 1'b0;
            15'b10000011_0101_010: DATA = 1'b0;
            15'b10000011_0101_011: DATA = 1'b1;
            15'b10000011_0101_100: DATA = 1'b1;
            15'b10000011_0101_101: DATA = 1'b0;
            15'b10000011_0101_110: DATA = 1'b0;
            15'b10000011_0101_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 3 Row 6
            15'b10000011_0110_000: DATA = 1'b0;
            15'b10000011_0110_001: DATA = 1'b0;
            15'b10000011_0110_010: DATA = 1'b0;
            15'b10000011_0110_011: DATA = 1'b0;
            15'b10000011_0110_100: DATA = 1'b1;
            15'b10000011_0110_101: DATA = 1'b1;
            15'b10000011_0110_110: DATA = 1'b0;
            15'b10000011_0110_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 3 Row 7
            15'b10000011_0111_000: DATA = 1'b0;
            15'b10000011_0111_001: DATA = 1'b0;
            15'b10000011_0111_010: DATA = 1'b0;
            15'b10000011_0111_011: DATA = 1'b0;
            15'b10000011_0111_100: DATA = 1'b0;
            15'b10000011_0111_101: DATA = 1'b1;
            15'b10000011_0111_110: DATA = 1'b1;
            15'b10000011_0111_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 3 Row 8
            15'b10000011_1000_000: DATA = 1'b0;
            15'b10000011_1000_001: DATA = 1'b0;
            15'b10000011_1000_010: DATA = 1'b0;
            15'b10000011_1000_011: DATA = 1'b0;
            15'b10000011_1000_100: DATA = 1'b0;
            15'b10000011_1000_101: DATA = 1'b0;
            15'b10000011_1000_110: DATA = 1'b1;
            15'b10000011_1000_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 3 Row 9
            15'b10000011_1001_000: DATA = 1'b0;
            15'b10000011_1001_001: DATA = 1'b0;
            15'b10000011_1001_010: DATA = 1'b0;
            15'b10000011_1001_011: DATA = 1'b0;
            15'b10000011_1001_100: DATA = 1'b0;
            15'b10000011_1001_101: DATA = 1'b0;
            15'b10000011_1001_110: DATA = 1'b1;
            15'b10000011_1001_111: DATA = 1'b1;
            // SINE+ ROW 0 COL 3 Row 10
            15'b10000011_1010_000: DATA = 1'b0;
            15'b10000011_1010_001: DATA = 1'b0;
            15'b10000011_1010_010: DATA = 1'b0;
            15'b10000011_1010_011: DATA = 1'b0;
            15'b10000011_1010_100: DATA = 1'b0;
            15'b10000011_1010_101: DATA = 1'b0;
            15'b10000011_1010_110: DATA = 1'b0;
            15'b10000011_1010_111: DATA = 1'b1;
            // SINE+ ROW 0 COL 3 Row 11
            15'b10000011_1011_000: DATA = 1'b0;
            15'b10000011_1011_001: DATA = 1'b0;
            15'b10000011_1011_010: DATA = 1'b0;
            15'b10000011_1011_011: DATA = 1'b0;
            15'b10000011_1011_100: DATA = 1'b0;
            15'b10000011_1011_101: DATA = 1'b0;
            15'b10000011_1011_110: DATA = 1'b0;
            15'b10000011_1011_111: DATA = 1'b1;
            // SINE+ ROW 0 COL 3 Row 12
            15'b10000011_1100_000: DATA = 1'b0;
            15'b10000011_1100_001: DATA = 1'b0;
            15'b10000011_1100_010: DATA = 1'b0;
            15'b10000011_1100_011: DATA = 1'b0;
            15'b10000011_1100_100: DATA = 1'b0;
            15'b10000011_1100_101: DATA = 1'b0;
            15'b10000011_1100_110: DATA = 1'b0;
            15'b10000011_1100_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 3 Row 13
            15'b10000011_1101_000: DATA = 1'b0;
            15'b10000011_1101_001: DATA = 1'b0;
            15'b10000011_1101_010: DATA = 1'b0;
            15'b10000011_1101_011: DATA = 1'b0;
            15'b10000011_1101_100: DATA = 1'b0;
            15'b10000011_1101_101: DATA = 1'b0;
            15'b10000011_1101_110: DATA = 1'b0;
            15'b10000011_1101_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 3 Row 14
            15'b10000011_1110_000: DATA = 1'b0;
            15'b10000011_1110_001: DATA = 1'b0;
            15'b10000011_1110_010: DATA = 1'b0;
            15'b10000011_1110_011: DATA = 1'b0;
            15'b10000011_1110_100: DATA = 1'b0;
            15'b10000011_1110_101: DATA = 1'b0;
            15'b10000011_1110_110: DATA = 1'b0;
            15'b10000011_1110_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 3 Row 15
            15'b10000011_1111_000: DATA = 1'b0;
            15'b10000011_1111_001: DATA = 1'b0;
            15'b10000011_1111_010: DATA = 1'b0;
            15'b10000011_1111_011: DATA = 1'b0;
            15'b10000011_1111_100: DATA = 1'b0;
            15'b10000011_1111_101: DATA = 1'b0;
            15'b10000011_1111_110: DATA = 1'b0;
            15'b10000011_1111_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 4 Row 0
            15'b10000100_0000_000: DATA = 1'b0;
            15'b10000100_0000_001: DATA = 1'b0;
            15'b10000100_0000_010: DATA = 1'b0;
            15'b10000100_0000_011: DATA = 1'b0;
            15'b10000100_0000_100: DATA = 1'b0;
            15'b10000100_0000_101: DATA = 1'b0;
            15'b10000100_0000_110: DATA = 1'b0;
            15'b10000100_0000_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 4 Row 1
            15'b10000100_0001_000: DATA = 1'b0;
            15'b10000100_0001_001: DATA = 1'b0;
            15'b10000100_0001_010: DATA = 1'b0;
            15'b10000100_0001_011: DATA = 1'b0;
            15'b10000100_0001_100: DATA = 1'b0;
            15'b10000100_0001_101: DATA = 1'b0;
            15'b10000100_0001_110: DATA = 1'b0;
            15'b10000100_0001_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 4 Row 2
            15'b10000100_0010_000: DATA = 1'b0;
            15'b10000100_0010_001: DATA = 1'b0;
            15'b10000100_0010_010: DATA = 1'b0;
            15'b10000100_0010_011: DATA = 1'b0;
            15'b10000100_0010_100: DATA = 1'b0;
            15'b10000100_0010_101: DATA = 1'b0;
            15'b10000100_0010_110: DATA = 1'b0;
            15'b10000100_0010_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 4 Row 3
            15'b10000100_0011_000: DATA = 1'b0;
            15'b10000100_0011_001: DATA = 1'b0;
            15'b10000100_0011_010: DATA = 1'b0;
            15'b10000100_0011_011: DATA = 1'b0;
            15'b10000100_0011_100: DATA = 1'b0;
            15'b10000100_0011_101: DATA = 1'b0;
            15'b10000100_0011_110: DATA = 1'b0;
            15'b10000100_0011_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 4 Row 4
            15'b10000100_0100_000: DATA = 1'b0;
            15'b10000100_0100_001: DATA = 1'b0;
            15'b10000100_0100_010: DATA = 1'b0;
            15'b10000100_0100_011: DATA = 1'b0;
            15'b10000100_0100_100: DATA = 1'b0;
            15'b10000100_0100_101: DATA = 1'b0;
            15'b10000100_0100_110: DATA = 1'b0;
            15'b10000100_0100_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 4 Row 5
            15'b10000100_0101_000: DATA = 1'b0;
            15'b10000100_0101_001: DATA = 1'b0;
            15'b10000100_0101_010: DATA = 1'b0;
            15'b10000100_0101_011: DATA = 1'b0;
            15'b10000100_0101_100: DATA = 1'b0;
            15'b10000100_0101_101: DATA = 1'b0;
            15'b10000100_0101_110: DATA = 1'b0;
            15'b10000100_0101_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 4 Row 6
            15'b10000100_0110_000: DATA = 1'b0;
            15'b10000100_0110_001: DATA = 1'b0;
            15'b10000100_0110_010: DATA = 1'b0;
            15'b10000100_0110_011: DATA = 1'b0;
            15'b10000100_0110_100: DATA = 1'b0;
            15'b10000100_0110_101: DATA = 1'b0;
            15'b10000100_0110_110: DATA = 1'b0;
            15'b10000100_0110_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 4 Row 7
            15'b10000100_0111_000: DATA = 1'b0;
            15'b10000100_0111_001: DATA = 1'b0;
            15'b10000100_0111_010: DATA = 1'b0;
            15'b10000100_0111_011: DATA = 1'b0;
            15'b10000100_0111_100: DATA = 1'b0;
            15'b10000100_0111_101: DATA = 1'b0;
            15'b10000100_0111_110: DATA = 1'b0;
            15'b10000100_0111_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 4 Row 8
            15'b10000100_1000_000: DATA = 1'b0;
            15'b10000100_1000_001: DATA = 1'b0;
            15'b10000100_1000_010: DATA = 1'b0;
            15'b10000100_1000_011: DATA = 1'b0;
            15'b10000100_1000_100: DATA = 1'b0;
            15'b10000100_1000_101: DATA = 1'b0;
            15'b10000100_1000_110: DATA = 1'b0;
            15'b10000100_1000_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 4 Row 9
            15'b10000100_1001_000: DATA = 1'b0;
            15'b10000100_1001_001: DATA = 1'b0;
            15'b10000100_1001_010: DATA = 1'b0;
            15'b10000100_1001_011: DATA = 1'b0;
            15'b10000100_1001_100: DATA = 1'b0;
            15'b10000100_1001_101: DATA = 1'b0;
            15'b10000100_1001_110: DATA = 1'b0;
            15'b10000100_1001_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 4 Row 10
            15'b10000100_1010_000: DATA = 1'b0;
            15'b10000100_1010_001: DATA = 1'b0;
            15'b10000100_1010_010: DATA = 1'b0;
            15'b10000100_1010_011: DATA = 1'b0;
            15'b10000100_1010_100: DATA = 1'b0;
            15'b10000100_1010_101: DATA = 1'b0;
            15'b10000100_1010_110: DATA = 1'b0;
            15'b10000100_1010_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 4 Row 11
            15'b10000100_1011_000: DATA = 1'b1;
            15'b10000100_1011_001: DATA = 1'b0;
            15'b10000100_1011_010: DATA = 1'b0;
            15'b10000100_1011_011: DATA = 1'b0;
            15'b10000100_1011_100: DATA = 1'b0;
            15'b10000100_1011_101: DATA = 1'b0;
            15'b10000100_1011_110: DATA = 1'b0;
            15'b10000100_1011_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 4 Row 12
            15'b10000100_1100_000: DATA = 1'b1;
            15'b10000100_1100_001: DATA = 1'b0;
            15'b10000100_1100_010: DATA = 1'b0;
            15'b10000100_1100_011: DATA = 1'b0;
            15'b10000100_1100_100: DATA = 1'b0;
            15'b10000100_1100_101: DATA = 1'b0;
            15'b10000100_1100_110: DATA = 1'b0;
            15'b10000100_1100_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 4 Row 13
            15'b10000100_1101_000: DATA = 1'b1;
            15'b10000100_1101_001: DATA = 1'b1;
            15'b10000100_1101_010: DATA = 1'b0;
            15'b10000100_1101_011: DATA = 1'b0;
            15'b10000100_1101_100: DATA = 1'b0;
            15'b10000100_1101_101: DATA = 1'b0;
            15'b10000100_1101_110: DATA = 1'b0;
            15'b10000100_1101_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 4 Row 14
            15'b10000100_1110_000: DATA = 1'b0;
            15'b10000100_1110_001: DATA = 1'b1;
            15'b10000100_1110_010: DATA = 1'b0;
            15'b10000100_1110_011: DATA = 1'b0;
            15'b10000100_1110_100: DATA = 1'b0;
            15'b10000100_1110_101: DATA = 1'b0;
            15'b10000100_1110_110: DATA = 1'b0;
            15'b10000100_1110_111: DATA = 1'b0;
            // SINE+ ROW 0 COL 4 Row 15
            15'b10000100_1111_000: DATA = 1'b0;
            15'b10000100_1111_001: DATA = 1'b1;
            15'b10000100_1111_010: DATA = 1'b1;
            15'b10000100_1111_011: DATA = 1'b0;
            15'b10000100_1111_100: DATA = 1'b0;
            15'b10000100_1111_101: DATA = 1'b0;
            15'b10000100_1111_110: DATA = 1'b0;
            15'b10000100_1111_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 0 Row 0
            15'b10000101_0000_000: DATA = 1'b0;
            15'b10000101_0000_001: DATA = 1'b0;
            15'b10000101_0000_010: DATA = 1'b0;
            15'b10000101_0000_011: DATA = 1'b0;
            15'b10000101_0000_100: DATA = 1'b0;
            15'b10000101_0000_101: DATA = 1'b1;
            15'b10000101_0000_110: DATA = 1'b0;
            15'b10000101_0000_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 0 Row 1
            15'b10000101_0001_000: DATA = 1'b0;
            15'b10000101_0001_001: DATA = 1'b0;
            15'b10000101_0001_010: DATA = 1'b0;
            15'b10000101_0001_011: DATA = 1'b0;
            15'b10000101_0001_100: DATA = 1'b1;
            15'b10000101_0001_101: DATA = 1'b1;
            15'b10000101_0001_110: DATA = 1'b0;
            15'b10000101_0001_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 0 Row 2
            15'b10000101_0010_000: DATA = 1'b0;
            15'b10000101_0010_001: DATA = 1'b0;
            15'b10000101_0010_010: DATA = 1'b0;
            15'b10000101_0010_011: DATA = 1'b0;
            15'b10000101_0010_100: DATA = 1'b1;
            15'b10000101_0010_101: DATA = 1'b0;
            15'b10000101_0010_110: DATA = 1'b0;
            15'b10000101_0010_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 0 Row 3
            15'b10000101_0011_000: DATA = 1'b0;
            15'b10000101_0011_001: DATA = 1'b0;
            15'b10000101_0011_010: DATA = 1'b0;
            15'b10000101_0011_011: DATA = 1'b1;
            15'b10000101_0011_100: DATA = 1'b1;
            15'b10000101_0011_101: DATA = 1'b0;
            15'b10000101_0011_110: DATA = 1'b0;
            15'b10000101_0011_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 0 Row 4
            15'b10000101_0100_000: DATA = 1'b0;
            15'b10000101_0100_001: DATA = 1'b0;
            15'b10000101_0100_010: DATA = 1'b0;
            15'b10000101_0100_011: DATA = 1'b1;
            15'b10000101_0100_100: DATA = 1'b0;
            15'b10000101_0100_101: DATA = 1'b0;
            15'b10000101_0100_110: DATA = 1'b0;
            15'b10000101_0100_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 0 Row 5
            15'b10000101_0101_000: DATA = 1'b0;
            15'b10000101_0101_001: DATA = 1'b0;
            15'b10000101_0101_010: DATA = 1'b0;
            15'b10000101_0101_011: DATA = 1'b1;
            15'b10000101_0101_100: DATA = 1'b0;
            15'b10000101_0101_101: DATA = 1'b0;
            15'b10000101_0101_110: DATA = 1'b0;
            15'b10000101_0101_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 0 Row 6
            15'b10000101_0110_000: DATA = 1'b0;
            15'b10000101_0110_001: DATA = 1'b0;
            15'b10000101_0110_010: DATA = 1'b1;
            15'b10000101_0110_011: DATA = 1'b1;
            15'b10000101_0110_100: DATA = 1'b0;
            15'b10000101_0110_101: DATA = 1'b0;
            15'b10000101_0110_110: DATA = 1'b0;
            15'b10000101_0110_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 0 Row 7
            15'b10000101_0111_000: DATA = 1'b0;
            15'b10000101_0111_001: DATA = 1'b0;
            15'b10000101_0111_010: DATA = 1'b1;
            15'b10000101_0111_011: DATA = 1'b0;
            15'b10000101_0111_100: DATA = 1'b0;
            15'b10000101_0111_101: DATA = 1'b0;
            15'b10000101_0111_110: DATA = 1'b0;
            15'b10000101_0111_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 0 Row 8
            15'b10000101_1000_000: DATA = 1'b0;
            15'b10000101_1000_001: DATA = 1'b0;
            15'b10000101_1000_010: DATA = 1'b1;
            15'b10000101_1000_011: DATA = 1'b0;
            15'b10000101_1000_100: DATA = 1'b0;
            15'b10000101_1000_101: DATA = 1'b0;
            15'b10000101_1000_110: DATA = 1'b0;
            15'b10000101_1000_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 0 Row 9
            15'b10000101_1001_000: DATA = 1'b0;
            15'b10000101_1001_001: DATA = 1'b1;
            15'b10000101_1001_010: DATA = 1'b1;
            15'b10000101_1001_011: DATA = 1'b0;
            15'b10000101_1001_100: DATA = 1'b0;
            15'b10000101_1001_101: DATA = 1'b0;
            15'b10000101_1001_110: DATA = 1'b0;
            15'b10000101_1001_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 0 Row 10
            15'b10000101_1010_000: DATA = 1'b0;
            15'b10000101_1010_001: DATA = 1'b1;
            15'b10000101_1010_010: DATA = 1'b0;
            15'b10000101_1010_011: DATA = 1'b0;
            15'b10000101_1010_100: DATA = 1'b0;
            15'b10000101_1010_101: DATA = 1'b0;
            15'b10000101_1010_110: DATA = 1'b0;
            15'b10000101_1010_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 0 Row 11
            15'b10000101_1011_000: DATA = 1'b0;
            15'b10000101_1011_001: DATA = 1'b1;
            15'b10000101_1011_010: DATA = 1'b0;
            15'b10000101_1011_011: DATA = 1'b0;
            15'b10000101_1011_100: DATA = 1'b0;
            15'b10000101_1011_101: DATA = 1'b0;
            15'b10000101_1011_110: DATA = 1'b0;
            15'b10000101_1011_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 0 Row 12
            15'b10000101_1100_000: DATA = 1'b1;
            15'b10000101_1100_001: DATA = 1'b1;
            15'b10000101_1100_010: DATA = 1'b0;
            15'b10000101_1100_011: DATA = 1'b0;
            15'b10000101_1100_100: DATA = 1'b0;
            15'b10000101_1100_101: DATA = 1'b0;
            15'b10000101_1100_110: DATA = 1'b0;
            15'b10000101_1100_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 0 Row 13
            15'b10000101_1101_000: DATA = 1'b1;
            15'b10000101_1101_001: DATA = 1'b0;
            15'b10000101_1101_010: DATA = 1'b0;
            15'b10000101_1101_011: DATA = 1'b0;
            15'b10000101_1101_100: DATA = 1'b0;
            15'b10000101_1101_101: DATA = 1'b0;
            15'b10000101_1101_110: DATA = 1'b0;
            15'b10000101_1101_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 0 Row 14
            15'b10000101_1110_000: DATA = 1'b1;
            15'b10000101_1110_001: DATA = 1'b0;
            15'b10000101_1110_010: DATA = 1'b0;
            15'b10000101_1110_011: DATA = 1'b0;
            15'b10000101_1110_100: DATA = 1'b0;
            15'b10000101_1110_101: DATA = 1'b0;
            15'b10000101_1110_110: DATA = 1'b0;
            15'b10000101_1110_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 0 Row 15
            15'b10000101_1111_000: DATA = 1'b1;
            15'b10000101_1111_001: DATA = 1'b0;
            15'b10000101_1111_010: DATA = 1'b0;
            15'b10000101_1111_011: DATA = 1'b0;
            15'b10000101_1111_100: DATA = 1'b0;
            15'b10000101_1111_101: DATA = 1'b0;
            15'b10000101_1111_110: DATA = 1'b0;
            15'b10000101_1111_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 1 Row 0
            15'b10000110_0000_000: DATA = 1'b0;
            15'b10000110_0000_001: DATA = 1'b0;
            15'b10000110_0000_010: DATA = 1'b0;
            15'b10000110_0000_011: DATA = 1'b0;
            15'b10000110_0000_100: DATA = 1'b0;
            15'b10000110_0000_101: DATA = 1'b0;
            15'b10000110_0000_110: DATA = 1'b0;
            15'b10000110_0000_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 1 Row 1
            15'b10000110_0001_000: DATA = 1'b0;
            15'b10000110_0001_001: DATA = 1'b0;
            15'b10000110_0001_010: DATA = 1'b0;
            15'b10000110_0001_011: DATA = 1'b0;
            15'b10000110_0001_100: DATA = 1'b0;
            15'b10000110_0001_101: DATA = 1'b0;
            15'b10000110_0001_110: DATA = 1'b0;
            15'b10000110_0001_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 1 Row 2
            15'b10000110_0010_000: DATA = 1'b0;
            15'b10000110_0010_001: DATA = 1'b0;
            15'b10000110_0010_010: DATA = 1'b0;
            15'b10000110_0010_011: DATA = 1'b0;
            15'b10000110_0010_100: DATA = 1'b0;
            15'b10000110_0010_101: DATA = 1'b0;
            15'b10000110_0010_110: DATA = 1'b0;
            15'b10000110_0010_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 1 Row 3
            15'b10000110_0011_000: DATA = 1'b0;
            15'b10000110_0011_001: DATA = 1'b0;
            15'b10000110_0011_010: DATA = 1'b0;
            15'b10000110_0011_011: DATA = 1'b0;
            15'b10000110_0011_100: DATA = 1'b0;
            15'b10000110_0011_101: DATA = 1'b0;
            15'b10000110_0011_110: DATA = 1'b0;
            15'b10000110_0011_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 1 Row 4
            15'b10000110_0100_000: DATA = 1'b0;
            15'b10000110_0100_001: DATA = 1'b0;
            15'b10000110_0100_010: DATA = 1'b0;
            15'b10000110_0100_011: DATA = 1'b0;
            15'b10000110_0100_100: DATA = 1'b0;
            15'b10000110_0100_101: DATA = 1'b0;
            15'b10000110_0100_110: DATA = 1'b0;
            15'b10000110_0100_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 1 Row 5
            15'b10000110_0101_000: DATA = 1'b0;
            15'b10000110_0101_001: DATA = 1'b0;
            15'b10000110_0101_010: DATA = 1'b0;
            15'b10000110_0101_011: DATA = 1'b0;
            15'b10000110_0101_100: DATA = 1'b0;
            15'b10000110_0101_101: DATA = 1'b0;
            15'b10000110_0101_110: DATA = 1'b0;
            15'b10000110_0101_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 1 Row 6
            15'b10000110_0110_000: DATA = 1'b0;
            15'b10000110_0110_001: DATA = 1'b0;
            15'b10000110_0110_010: DATA = 1'b0;
            15'b10000110_0110_011: DATA = 1'b0;
            15'b10000110_0110_100: DATA = 1'b0;
            15'b10000110_0110_101: DATA = 1'b0;
            15'b10000110_0110_110: DATA = 1'b0;
            15'b10000110_0110_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 1 Row 7
            15'b10000110_0111_000: DATA = 1'b0;
            15'b10000110_0111_001: DATA = 1'b0;
            15'b10000110_0111_010: DATA = 1'b0;
            15'b10000110_0111_011: DATA = 1'b0;
            15'b10000110_0111_100: DATA = 1'b0;
            15'b10000110_0111_101: DATA = 1'b0;
            15'b10000110_0111_110: DATA = 1'b0;
            15'b10000110_0111_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 1 Row 8
            15'b10000110_1000_000: DATA = 1'b0;
            15'b10000110_1000_001: DATA = 1'b0;
            15'b10000110_1000_010: DATA = 1'b0;
            15'b10000110_1000_011: DATA = 1'b0;
            15'b10000110_1000_100: DATA = 1'b0;
            15'b10000110_1000_101: DATA = 1'b0;
            15'b10000110_1000_110: DATA = 1'b0;
            15'b10000110_1000_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 1 Row 9
            15'b10000110_1001_000: DATA = 1'b0;
            15'b10000110_1001_001: DATA = 1'b0;
            15'b10000110_1001_010: DATA = 1'b0;
            15'b10000110_1001_011: DATA = 1'b0;
            15'b10000110_1001_100: DATA = 1'b0;
            15'b10000110_1001_101: DATA = 1'b0;
            15'b10000110_1001_110: DATA = 1'b0;
            15'b10000110_1001_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 1 Row 10
            15'b10000110_1010_000: DATA = 1'b0;
            15'b10000110_1010_001: DATA = 1'b0;
            15'b10000110_1010_010: DATA = 1'b0;
            15'b10000110_1010_011: DATA = 1'b0;
            15'b10000110_1010_100: DATA = 1'b0;
            15'b10000110_1010_101: DATA = 1'b0;
            15'b10000110_1010_110: DATA = 1'b0;
            15'b10000110_1010_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 1 Row 11
            15'b10000110_1011_000: DATA = 1'b0;
            15'b10000110_1011_001: DATA = 1'b0;
            15'b10000110_1011_010: DATA = 1'b0;
            15'b10000110_1011_011: DATA = 1'b0;
            15'b10000110_1011_100: DATA = 1'b0;
            15'b10000110_1011_101: DATA = 1'b0;
            15'b10000110_1011_110: DATA = 1'b0;
            15'b10000110_1011_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 1 Row 12
            15'b10000110_1100_000: DATA = 1'b0;
            15'b10000110_1100_001: DATA = 1'b0;
            15'b10000110_1100_010: DATA = 1'b0;
            15'b10000110_1100_011: DATA = 1'b0;
            15'b10000110_1100_100: DATA = 1'b0;
            15'b10000110_1100_101: DATA = 1'b0;
            15'b10000110_1100_110: DATA = 1'b0;
            15'b10000110_1100_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 1 Row 13
            15'b10000110_1101_000: DATA = 1'b0;
            15'b10000110_1101_001: DATA = 1'b0;
            15'b10000110_1101_010: DATA = 1'b0;
            15'b10000110_1101_011: DATA = 1'b0;
            15'b10000110_1101_100: DATA = 1'b0;
            15'b10000110_1101_101: DATA = 1'b0;
            15'b10000110_1101_110: DATA = 1'b0;
            15'b10000110_1101_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 1 Row 14
            15'b10000110_1110_000: DATA = 1'b0;
            15'b10000110_1110_001: DATA = 1'b0;
            15'b10000110_1110_010: DATA = 1'b0;
            15'b10000110_1110_011: DATA = 1'b0;
            15'b10000110_1110_100: DATA = 1'b0;
            15'b10000110_1110_101: DATA = 1'b0;
            15'b10000110_1110_110: DATA = 1'b0;
            15'b10000110_1110_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 1 Row 15
            15'b10000110_1111_000: DATA = 1'b0;
            15'b10000110_1111_001: DATA = 1'b0;
            15'b10000110_1111_010: DATA = 1'b0;
            15'b10000110_1111_011: DATA = 1'b0;
            15'b10000110_1111_100: DATA = 1'b0;
            15'b10000110_1111_101: DATA = 1'b0;
            15'b10000110_1111_110: DATA = 1'b0;
            15'b10000110_1111_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 2 Row 0
            15'b10000111_0000_000: DATA = 1'b0;
            15'b10000111_0000_001: DATA = 1'b0;
            15'b10000111_0000_010: DATA = 1'b0;
            15'b10000111_0000_011: DATA = 1'b0;
            15'b10000111_0000_100: DATA = 1'b0;
            15'b10000111_0000_101: DATA = 1'b0;
            15'b10000111_0000_110: DATA = 1'b0;
            15'b10000111_0000_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 2 Row 1
            15'b10000111_0001_000: DATA = 1'b0;
            15'b10000111_0001_001: DATA = 1'b0;
            15'b10000111_0001_010: DATA = 1'b0;
            15'b10000111_0001_011: DATA = 1'b0;
            15'b10000111_0001_100: DATA = 1'b0;
            15'b10000111_0001_101: DATA = 1'b0;
            15'b10000111_0001_110: DATA = 1'b0;
            15'b10000111_0001_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 2 Row 2
            15'b10000111_0010_000: DATA = 1'b0;
            15'b10000111_0010_001: DATA = 1'b0;
            15'b10000111_0010_010: DATA = 1'b0;
            15'b10000111_0010_011: DATA = 1'b0;
            15'b10000111_0010_100: DATA = 1'b0;
            15'b10000111_0010_101: DATA = 1'b0;
            15'b10000111_0010_110: DATA = 1'b0;
            15'b10000111_0010_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 2 Row 3
            15'b10000111_0011_000: DATA = 1'b0;
            15'b10000111_0011_001: DATA = 1'b0;
            15'b10000111_0011_010: DATA = 1'b0;
            15'b10000111_0011_011: DATA = 1'b0;
            15'b10000111_0011_100: DATA = 1'b0;
            15'b10000111_0011_101: DATA = 1'b0;
            15'b10000111_0011_110: DATA = 1'b0;
            15'b10000111_0011_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 2 Row 4
            15'b10000111_0100_000: DATA = 1'b0;
            15'b10000111_0100_001: DATA = 1'b0;
            15'b10000111_0100_010: DATA = 1'b0;
            15'b10000111_0100_011: DATA = 1'b0;
            15'b10000111_0100_100: DATA = 1'b0;
            15'b10000111_0100_101: DATA = 1'b0;
            15'b10000111_0100_110: DATA = 1'b0;
            15'b10000111_0100_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 2 Row 5
            15'b10000111_0101_000: DATA = 1'b0;
            15'b10000111_0101_001: DATA = 1'b0;
            15'b10000111_0101_010: DATA = 1'b0;
            15'b10000111_0101_011: DATA = 1'b0;
            15'b10000111_0101_100: DATA = 1'b0;
            15'b10000111_0101_101: DATA = 1'b0;
            15'b10000111_0101_110: DATA = 1'b0;
            15'b10000111_0101_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 2 Row 6
            15'b10000111_0110_000: DATA = 1'b0;
            15'b10000111_0110_001: DATA = 1'b0;
            15'b10000111_0110_010: DATA = 1'b0;
            15'b10000111_0110_011: DATA = 1'b0;
            15'b10000111_0110_100: DATA = 1'b0;
            15'b10000111_0110_101: DATA = 1'b0;
            15'b10000111_0110_110: DATA = 1'b0;
            15'b10000111_0110_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 2 Row 7
            15'b10000111_0111_000: DATA = 1'b0;
            15'b10000111_0111_001: DATA = 1'b0;
            15'b10000111_0111_010: DATA = 1'b0;
            15'b10000111_0111_011: DATA = 1'b0;
            15'b10000111_0111_100: DATA = 1'b0;
            15'b10000111_0111_101: DATA = 1'b0;
            15'b10000111_0111_110: DATA = 1'b0;
            15'b10000111_0111_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 2 Row 8
            15'b10000111_1000_000: DATA = 1'b0;
            15'b10000111_1000_001: DATA = 1'b0;
            15'b10000111_1000_010: DATA = 1'b0;
            15'b10000111_1000_011: DATA = 1'b0;
            15'b10000111_1000_100: DATA = 1'b0;
            15'b10000111_1000_101: DATA = 1'b0;
            15'b10000111_1000_110: DATA = 1'b0;
            15'b10000111_1000_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 2 Row 9
            15'b10000111_1001_000: DATA = 1'b0;
            15'b10000111_1001_001: DATA = 1'b0;
            15'b10000111_1001_010: DATA = 1'b0;
            15'b10000111_1001_011: DATA = 1'b0;
            15'b10000111_1001_100: DATA = 1'b0;
            15'b10000111_1001_101: DATA = 1'b0;
            15'b10000111_1001_110: DATA = 1'b0;
            15'b10000111_1001_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 2 Row 10
            15'b10000111_1010_000: DATA = 1'b0;
            15'b10000111_1010_001: DATA = 1'b0;
            15'b10000111_1010_010: DATA = 1'b0;
            15'b10000111_1010_011: DATA = 1'b0;
            15'b10000111_1010_100: DATA = 1'b0;
            15'b10000111_1010_101: DATA = 1'b0;
            15'b10000111_1010_110: DATA = 1'b0;
            15'b10000111_1010_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 2 Row 11
            15'b10000111_1011_000: DATA = 1'b0;
            15'b10000111_1011_001: DATA = 1'b0;
            15'b10000111_1011_010: DATA = 1'b0;
            15'b10000111_1011_011: DATA = 1'b0;
            15'b10000111_1011_100: DATA = 1'b0;
            15'b10000111_1011_101: DATA = 1'b0;
            15'b10000111_1011_110: DATA = 1'b0;
            15'b10000111_1011_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 2 Row 12
            15'b10000111_1100_000: DATA = 1'b0;
            15'b10000111_1100_001: DATA = 1'b0;
            15'b10000111_1100_010: DATA = 1'b0;
            15'b10000111_1100_011: DATA = 1'b0;
            15'b10000111_1100_100: DATA = 1'b0;
            15'b10000111_1100_101: DATA = 1'b0;
            15'b10000111_1100_110: DATA = 1'b0;
            15'b10000111_1100_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 2 Row 13
            15'b10000111_1101_000: DATA = 1'b0;
            15'b10000111_1101_001: DATA = 1'b0;
            15'b10000111_1101_010: DATA = 1'b0;
            15'b10000111_1101_011: DATA = 1'b0;
            15'b10000111_1101_100: DATA = 1'b0;
            15'b10000111_1101_101: DATA = 1'b0;
            15'b10000111_1101_110: DATA = 1'b0;
            15'b10000111_1101_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 2 Row 14
            15'b10000111_1110_000: DATA = 1'b0;
            15'b10000111_1110_001: DATA = 1'b0;
            15'b10000111_1110_010: DATA = 1'b0;
            15'b10000111_1110_011: DATA = 1'b0;
            15'b10000111_1110_100: DATA = 1'b0;
            15'b10000111_1110_101: DATA = 1'b0;
            15'b10000111_1110_110: DATA = 1'b0;
            15'b10000111_1110_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 2 Row 15
            15'b10000111_1111_000: DATA = 1'b0;
            15'b10000111_1111_001: DATA = 1'b0;
            15'b10000111_1111_010: DATA = 1'b0;
            15'b10000111_1111_011: DATA = 1'b0;
            15'b10000111_1111_100: DATA = 1'b0;
            15'b10000111_1111_101: DATA = 1'b0;
            15'b10000111_1111_110: DATA = 1'b0;
            15'b10000111_1111_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 3 Row 0
            15'b10001000_0000_000: DATA = 1'b0;
            15'b10001000_0000_001: DATA = 1'b0;
            15'b10001000_0000_010: DATA = 1'b0;
            15'b10001000_0000_011: DATA = 1'b0;
            15'b10001000_0000_100: DATA = 1'b0;
            15'b10001000_0000_101: DATA = 1'b0;
            15'b10001000_0000_110: DATA = 1'b0;
            15'b10001000_0000_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 3 Row 1
            15'b10001000_0001_000: DATA = 1'b0;
            15'b10001000_0001_001: DATA = 1'b0;
            15'b10001000_0001_010: DATA = 1'b0;
            15'b10001000_0001_011: DATA = 1'b0;
            15'b10001000_0001_100: DATA = 1'b0;
            15'b10001000_0001_101: DATA = 1'b0;
            15'b10001000_0001_110: DATA = 1'b0;
            15'b10001000_0001_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 3 Row 2
            15'b10001000_0010_000: DATA = 1'b0;
            15'b10001000_0010_001: DATA = 1'b0;
            15'b10001000_0010_010: DATA = 1'b0;
            15'b10001000_0010_011: DATA = 1'b0;
            15'b10001000_0010_100: DATA = 1'b0;
            15'b10001000_0010_101: DATA = 1'b0;
            15'b10001000_0010_110: DATA = 1'b0;
            15'b10001000_0010_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 3 Row 3
            15'b10001000_0011_000: DATA = 1'b0;
            15'b10001000_0011_001: DATA = 1'b0;
            15'b10001000_0011_010: DATA = 1'b0;
            15'b10001000_0011_011: DATA = 1'b0;
            15'b10001000_0011_100: DATA = 1'b0;
            15'b10001000_0011_101: DATA = 1'b0;
            15'b10001000_0011_110: DATA = 1'b0;
            15'b10001000_0011_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 3 Row 4
            15'b10001000_0100_000: DATA = 1'b0;
            15'b10001000_0100_001: DATA = 1'b0;
            15'b10001000_0100_010: DATA = 1'b0;
            15'b10001000_0100_011: DATA = 1'b0;
            15'b10001000_0100_100: DATA = 1'b0;
            15'b10001000_0100_101: DATA = 1'b0;
            15'b10001000_0100_110: DATA = 1'b0;
            15'b10001000_0100_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 3 Row 5
            15'b10001000_0101_000: DATA = 1'b0;
            15'b10001000_0101_001: DATA = 1'b0;
            15'b10001000_0101_010: DATA = 1'b0;
            15'b10001000_0101_011: DATA = 1'b0;
            15'b10001000_0101_100: DATA = 1'b0;
            15'b10001000_0101_101: DATA = 1'b0;
            15'b10001000_0101_110: DATA = 1'b0;
            15'b10001000_0101_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 3 Row 6
            15'b10001000_0110_000: DATA = 1'b0;
            15'b10001000_0110_001: DATA = 1'b0;
            15'b10001000_0110_010: DATA = 1'b0;
            15'b10001000_0110_011: DATA = 1'b0;
            15'b10001000_0110_100: DATA = 1'b0;
            15'b10001000_0110_101: DATA = 1'b0;
            15'b10001000_0110_110: DATA = 1'b0;
            15'b10001000_0110_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 3 Row 7
            15'b10001000_0111_000: DATA = 1'b0;
            15'b10001000_0111_001: DATA = 1'b0;
            15'b10001000_0111_010: DATA = 1'b0;
            15'b10001000_0111_011: DATA = 1'b0;
            15'b10001000_0111_100: DATA = 1'b0;
            15'b10001000_0111_101: DATA = 1'b0;
            15'b10001000_0111_110: DATA = 1'b0;
            15'b10001000_0111_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 3 Row 8
            15'b10001000_1000_000: DATA = 1'b0;
            15'b10001000_1000_001: DATA = 1'b0;
            15'b10001000_1000_010: DATA = 1'b0;
            15'b10001000_1000_011: DATA = 1'b0;
            15'b10001000_1000_100: DATA = 1'b0;
            15'b10001000_1000_101: DATA = 1'b0;
            15'b10001000_1000_110: DATA = 1'b0;
            15'b10001000_1000_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 3 Row 9
            15'b10001000_1001_000: DATA = 1'b0;
            15'b10001000_1001_001: DATA = 1'b0;
            15'b10001000_1001_010: DATA = 1'b0;
            15'b10001000_1001_011: DATA = 1'b0;
            15'b10001000_1001_100: DATA = 1'b0;
            15'b10001000_1001_101: DATA = 1'b0;
            15'b10001000_1001_110: DATA = 1'b0;
            15'b10001000_1001_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 3 Row 10
            15'b10001000_1010_000: DATA = 1'b0;
            15'b10001000_1010_001: DATA = 1'b0;
            15'b10001000_1010_010: DATA = 1'b0;
            15'b10001000_1010_011: DATA = 1'b0;
            15'b10001000_1010_100: DATA = 1'b0;
            15'b10001000_1010_101: DATA = 1'b0;
            15'b10001000_1010_110: DATA = 1'b0;
            15'b10001000_1010_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 3 Row 11
            15'b10001000_1011_000: DATA = 1'b0;
            15'b10001000_1011_001: DATA = 1'b0;
            15'b10001000_1011_010: DATA = 1'b0;
            15'b10001000_1011_011: DATA = 1'b0;
            15'b10001000_1011_100: DATA = 1'b0;
            15'b10001000_1011_101: DATA = 1'b0;
            15'b10001000_1011_110: DATA = 1'b0;
            15'b10001000_1011_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 3 Row 12
            15'b10001000_1100_000: DATA = 1'b0;
            15'b10001000_1100_001: DATA = 1'b0;
            15'b10001000_1100_010: DATA = 1'b0;
            15'b10001000_1100_011: DATA = 1'b0;
            15'b10001000_1100_100: DATA = 1'b0;
            15'b10001000_1100_101: DATA = 1'b0;
            15'b10001000_1100_110: DATA = 1'b0;
            15'b10001000_1100_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 3 Row 13
            15'b10001000_1101_000: DATA = 1'b0;
            15'b10001000_1101_001: DATA = 1'b0;
            15'b10001000_1101_010: DATA = 1'b0;
            15'b10001000_1101_011: DATA = 1'b0;
            15'b10001000_1101_100: DATA = 1'b0;
            15'b10001000_1101_101: DATA = 1'b0;
            15'b10001000_1101_110: DATA = 1'b0;
            15'b10001000_1101_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 3 Row 14
            15'b10001000_1110_000: DATA = 1'b0;
            15'b10001000_1110_001: DATA = 1'b0;
            15'b10001000_1110_010: DATA = 1'b0;
            15'b10001000_1110_011: DATA = 1'b0;
            15'b10001000_1110_100: DATA = 1'b0;
            15'b10001000_1110_101: DATA = 1'b0;
            15'b10001000_1110_110: DATA = 1'b0;
            15'b10001000_1110_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 3 Row 15
            15'b10001000_1111_000: DATA = 1'b0;
            15'b10001000_1111_001: DATA = 1'b0;
            15'b10001000_1111_010: DATA = 1'b0;
            15'b10001000_1111_011: DATA = 1'b0;
            15'b10001000_1111_100: DATA = 1'b0;
            15'b10001000_1111_101: DATA = 1'b0;
            15'b10001000_1111_110: DATA = 1'b0;
            15'b10001000_1111_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 4 Row 0
            15'b10001001_0000_000: DATA = 1'b0;
            15'b10001001_0000_001: DATA = 1'b0;
            15'b10001001_0000_010: DATA = 1'b1;
            15'b10001001_0000_011: DATA = 1'b0;
            15'b10001001_0000_100: DATA = 1'b0;
            15'b10001001_0000_101: DATA = 1'b0;
            15'b10001001_0000_110: DATA = 1'b0;
            15'b10001001_0000_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 4 Row 1
            15'b10001001_0001_000: DATA = 1'b0;
            15'b10001001_0001_001: DATA = 1'b0;
            15'b10001001_0001_010: DATA = 1'b1;
            15'b10001001_0001_011: DATA = 1'b1;
            15'b10001001_0001_100: DATA = 1'b0;
            15'b10001001_0001_101: DATA = 1'b0;
            15'b10001001_0001_110: DATA = 1'b0;
            15'b10001001_0001_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 4 Row 2
            15'b10001001_0010_000: DATA = 1'b0;
            15'b10001001_0010_001: DATA = 1'b0;
            15'b10001001_0010_010: DATA = 1'b0;
            15'b10001001_0010_011: DATA = 1'b1;
            15'b10001001_0010_100: DATA = 1'b0;
            15'b10001001_0010_101: DATA = 1'b0;
            15'b10001001_0010_110: DATA = 1'b0;
            15'b10001001_0010_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 4 Row 3
            15'b10001001_0011_000: DATA = 1'b0;
            15'b10001001_0011_001: DATA = 1'b0;
            15'b10001001_0011_010: DATA = 1'b0;
            15'b10001001_0011_011: DATA = 1'b1;
            15'b10001001_0011_100: DATA = 1'b1;
            15'b10001001_0011_101: DATA = 1'b0;
            15'b10001001_0011_110: DATA = 1'b0;
            15'b10001001_0011_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 4 Row 4
            15'b10001001_0100_000: DATA = 1'b0;
            15'b10001001_0100_001: DATA = 1'b0;
            15'b10001001_0100_010: DATA = 1'b0;
            15'b10001001_0100_011: DATA = 1'b0;
            15'b10001001_0100_100: DATA = 1'b1;
            15'b10001001_0100_101: DATA = 1'b0;
            15'b10001001_0100_110: DATA = 1'b0;
            15'b10001001_0100_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 4 Row 5
            15'b10001001_0101_000: DATA = 1'b0;
            15'b10001001_0101_001: DATA = 1'b0;
            15'b10001001_0101_010: DATA = 1'b0;
            15'b10001001_0101_011: DATA = 1'b0;
            15'b10001001_0101_100: DATA = 1'b1;
            15'b10001001_0101_101: DATA = 1'b0;
            15'b10001001_0101_110: DATA = 1'b0;
            15'b10001001_0101_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 4 Row 6
            15'b10001001_0110_000: DATA = 1'b0;
            15'b10001001_0110_001: DATA = 1'b0;
            15'b10001001_0110_010: DATA = 1'b0;
            15'b10001001_0110_011: DATA = 1'b0;
            15'b10001001_0110_100: DATA = 1'b1;
            15'b10001001_0110_101: DATA = 1'b1;
            15'b10001001_0110_110: DATA = 1'b0;
            15'b10001001_0110_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 4 Row 7
            15'b10001001_0111_000: DATA = 1'b0;
            15'b10001001_0111_001: DATA = 1'b0;
            15'b10001001_0111_010: DATA = 1'b0;
            15'b10001001_0111_011: DATA = 1'b0;
            15'b10001001_0111_100: DATA = 1'b0;
            15'b10001001_0111_101: DATA = 1'b1;
            15'b10001001_0111_110: DATA = 1'b0;
            15'b10001001_0111_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 4 Row 8
            15'b10001001_1000_000: DATA = 1'b0;
            15'b10001001_1000_001: DATA = 1'b0;
            15'b10001001_1000_010: DATA = 1'b0;
            15'b10001001_1000_011: DATA = 1'b0;
            15'b10001001_1000_100: DATA = 1'b0;
            15'b10001001_1000_101: DATA = 1'b1;
            15'b10001001_1000_110: DATA = 1'b0;
            15'b10001001_1000_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 4 Row 9
            15'b10001001_1001_000: DATA = 1'b0;
            15'b10001001_1001_001: DATA = 1'b0;
            15'b10001001_1001_010: DATA = 1'b0;
            15'b10001001_1001_011: DATA = 1'b0;
            15'b10001001_1001_100: DATA = 1'b0;
            15'b10001001_1001_101: DATA = 1'b1;
            15'b10001001_1001_110: DATA = 1'b1;
            15'b10001001_1001_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 4 Row 10
            15'b10001001_1010_000: DATA = 1'b0;
            15'b10001001_1010_001: DATA = 1'b0;
            15'b10001001_1010_010: DATA = 1'b0;
            15'b10001001_1010_011: DATA = 1'b0;
            15'b10001001_1010_100: DATA = 1'b0;
            15'b10001001_1010_101: DATA = 1'b0;
            15'b10001001_1010_110: DATA = 1'b1;
            15'b10001001_1010_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 4 Row 11
            15'b10001001_1011_000: DATA = 1'b0;
            15'b10001001_1011_001: DATA = 1'b0;
            15'b10001001_1011_010: DATA = 1'b0;
            15'b10001001_1011_011: DATA = 1'b0;
            15'b10001001_1011_100: DATA = 1'b0;
            15'b10001001_1011_101: DATA = 1'b0;
            15'b10001001_1011_110: DATA = 1'b1;
            15'b10001001_1011_111: DATA = 1'b0;
            // SINE+ ROW 1 COL 4 Row 12
            15'b10001001_1100_000: DATA = 1'b0;
            15'b10001001_1100_001: DATA = 1'b0;
            15'b10001001_1100_010: DATA = 1'b0;
            15'b10001001_1100_011: DATA = 1'b0;
            15'b10001001_1100_100: DATA = 1'b0;
            15'b10001001_1100_101: DATA = 1'b0;
            15'b10001001_1100_110: DATA = 1'b1;
            15'b10001001_1100_111: DATA = 1'b1;
            // SINE+ ROW 1 COL 4 Row 13
            15'b10001001_1101_000: DATA = 1'b0;
            15'b10001001_1101_001: DATA = 1'b0;
            15'b10001001_1101_010: DATA = 1'b0;
            15'b10001001_1101_011: DATA = 1'b0;
            15'b10001001_1101_100: DATA = 1'b0;
            15'b10001001_1101_101: DATA = 1'b0;
            15'b10001001_1101_110: DATA = 1'b0;
            15'b10001001_1101_111: DATA = 1'b1;
            // SINE+ ROW 1 COL 4 Row 14
            15'b10001001_1110_000: DATA = 1'b0;
            15'b10001001_1110_001: DATA = 1'b0;
            15'b10001001_1110_010: DATA = 1'b0;
            15'b10001001_1110_011: DATA = 1'b0;
            15'b10001001_1110_100: DATA = 1'b0;
            15'b10001001_1110_101: DATA = 1'b0;
            15'b10001001_1110_110: DATA = 1'b0;
            15'b10001001_1110_111: DATA = 1'b1;
            // SINE+ ROW 1 COL 4 Row 15
            15'b10001001_1111_000: DATA = 1'b0;
            15'b10001001_1111_001: DATA = 1'b0;
            15'b10001001_1111_010: DATA = 1'b0;
            15'b10001001_1111_011: DATA = 1'b0;
            15'b10001001_1111_100: DATA = 1'b0;
            15'b10001001_1111_101: DATA = 1'b0;
            15'b10001001_1111_110: DATA = 1'b0;
            15'b10001001_1111_111: DATA = 1'b1;
            // SINE- ROW 0 COL 0 Row 0
            15'b10001010_0000_000: DATA = 1'b1;
            15'b10001010_0000_001: DATA = 1'b0;
            15'b10001010_0000_010: DATA = 1'b0;
            15'b10001010_0000_011: DATA = 1'b0;
            15'b10001010_0000_100: DATA = 1'b0;
            15'b10001010_0000_101: DATA = 1'b0;
            15'b10001010_0000_110: DATA = 1'b0;
            15'b10001010_0000_111: DATA = 1'b0;
            // SINE- ROW 0 COL 0 Row 1
            15'b10001010_0001_000: DATA = 1'b1;
            15'b10001010_0001_001: DATA = 1'b0;
            15'b10001010_0001_010: DATA = 1'b0;
            15'b10001010_0001_011: DATA = 1'b0;
            15'b10001010_0001_100: DATA = 1'b0;
            15'b10001010_0001_101: DATA = 1'b0;
            15'b10001010_0001_110: DATA = 1'b0;
            15'b10001010_0001_111: DATA = 1'b0;
            // SINE- ROW 0 COL 0 Row 2
            15'b10001010_0010_000: DATA = 1'b1;
            15'b10001010_0010_001: DATA = 1'b0;
            15'b10001010_0010_010: DATA = 1'b0;
            15'b10001010_0010_011: DATA = 1'b0;
            15'b10001010_0010_100: DATA = 1'b0;
            15'b10001010_0010_101: DATA = 1'b0;
            15'b10001010_0010_110: DATA = 1'b0;
            15'b10001010_0010_111: DATA = 1'b0;
            // SINE- ROW 0 COL 0 Row 3
            15'b10001010_0011_000: DATA = 1'b1;
            15'b10001010_0011_001: DATA = 1'b1;
            15'b10001010_0011_010: DATA = 1'b0;
            15'b10001010_0011_011: DATA = 1'b0;
            15'b10001010_0011_100: DATA = 1'b0;
            15'b10001010_0011_101: DATA = 1'b0;
            15'b10001010_0011_110: DATA = 1'b0;
            15'b10001010_0011_111: DATA = 1'b0;
            // SINE- ROW 0 COL 0 Row 4
            15'b10001010_0100_000: DATA = 1'b0;
            15'b10001010_0100_001: DATA = 1'b1;
            15'b10001010_0100_010: DATA = 1'b0;
            15'b10001010_0100_011: DATA = 1'b0;
            15'b10001010_0100_100: DATA = 1'b0;
            15'b10001010_0100_101: DATA = 1'b0;
            15'b10001010_0100_110: DATA = 1'b0;
            15'b10001010_0100_111: DATA = 1'b0;
            // SINE- ROW 0 COL 0 Row 5
            15'b10001010_0101_000: DATA = 1'b0;
            15'b10001010_0101_001: DATA = 1'b1;
            15'b10001010_0101_010: DATA = 1'b0;
            15'b10001010_0101_011: DATA = 1'b0;
            15'b10001010_0101_100: DATA = 1'b0;
            15'b10001010_0101_101: DATA = 1'b0;
            15'b10001010_0101_110: DATA = 1'b0;
            15'b10001010_0101_111: DATA = 1'b0;
            // SINE- ROW 0 COL 0 Row 6
            15'b10001010_0110_000: DATA = 1'b0;
            15'b10001010_0110_001: DATA = 1'b1;
            15'b10001010_0110_010: DATA = 1'b1;
            15'b10001010_0110_011: DATA = 1'b0;
            15'b10001010_0110_100: DATA = 1'b0;
            15'b10001010_0110_101: DATA = 1'b0;
            15'b10001010_0110_110: DATA = 1'b0;
            15'b10001010_0110_111: DATA = 1'b0;
            // SINE- ROW 0 COL 0 Row 7
            15'b10001010_0111_000: DATA = 1'b0;
            15'b10001010_0111_001: DATA = 1'b0;
            15'b10001010_0111_010: DATA = 1'b1;
            15'b10001010_0111_011: DATA = 1'b0;
            15'b10001010_0111_100: DATA = 1'b0;
            15'b10001010_0111_101: DATA = 1'b0;
            15'b10001010_0111_110: DATA = 1'b0;
            15'b10001010_0111_111: DATA = 1'b0;
            // SINE- ROW 0 COL 0 Row 8
            15'b10001010_1000_000: DATA = 1'b0;
            15'b10001010_1000_001: DATA = 1'b0;
            15'b10001010_1000_010: DATA = 1'b1;
            15'b10001010_1000_011: DATA = 1'b0;
            15'b10001010_1000_100: DATA = 1'b0;
            15'b10001010_1000_101: DATA = 1'b0;
            15'b10001010_1000_110: DATA = 1'b0;
            15'b10001010_1000_111: DATA = 1'b0;
            // SINE- ROW 0 COL 0 Row 9
            15'b10001010_1001_000: DATA = 1'b0;
            15'b10001010_1001_001: DATA = 1'b0;
            15'b10001010_1001_010: DATA = 1'b1;
            15'b10001010_1001_011: DATA = 1'b1;
            15'b10001010_1001_100: DATA = 1'b0;
            15'b10001010_1001_101: DATA = 1'b0;
            15'b10001010_1001_110: DATA = 1'b0;
            15'b10001010_1001_111: DATA = 1'b0;
            // SINE- ROW 0 COL 0 Row 10
            15'b10001010_1010_000: DATA = 1'b0;
            15'b10001010_1010_001: DATA = 1'b0;
            15'b10001010_1010_010: DATA = 1'b0;
            15'b10001010_1010_011: DATA = 1'b1;
            15'b10001010_1010_100: DATA = 1'b0;
            15'b10001010_1010_101: DATA = 1'b0;
            15'b10001010_1010_110: DATA = 1'b0;
            15'b10001010_1010_111: DATA = 1'b0;
            // SINE- ROW 0 COL 0 Row 11
            15'b10001010_1011_000: DATA = 1'b0;
            15'b10001010_1011_001: DATA = 1'b0;
            15'b10001010_1011_010: DATA = 1'b0;
            15'b10001010_1011_011: DATA = 1'b1;
            15'b10001010_1011_100: DATA = 1'b0;
            15'b10001010_1011_101: DATA = 1'b0;
            15'b10001010_1011_110: DATA = 1'b0;
            15'b10001010_1011_111: DATA = 1'b0;
            // SINE- ROW 0 COL 0 Row 12
            15'b10001010_1100_000: DATA = 1'b0;
            15'b10001010_1100_001: DATA = 1'b0;
            15'b10001010_1100_010: DATA = 1'b0;
            15'b10001010_1100_011: DATA = 1'b1;
            15'b10001010_1100_100: DATA = 1'b1;
            15'b10001010_1100_101: DATA = 1'b0;
            15'b10001010_1100_110: DATA = 1'b0;
            15'b10001010_1100_111: DATA = 1'b0;
            // SINE- ROW 0 COL 0 Row 13
            15'b10001010_1101_000: DATA = 1'b0;
            15'b10001010_1101_001: DATA = 1'b0;
            15'b10001010_1101_010: DATA = 1'b0;
            15'b10001010_1101_011: DATA = 1'b0;
            15'b10001010_1101_100: DATA = 1'b1;
            15'b10001010_1101_101: DATA = 1'b0;
            15'b10001010_1101_110: DATA = 1'b0;
            15'b10001010_1101_111: DATA = 1'b0;
            // SINE- ROW 0 COL 0 Row 14
            15'b10001010_1110_000: DATA = 1'b0;
            15'b10001010_1110_001: DATA = 1'b0;
            15'b10001010_1110_010: DATA = 1'b0;
            15'b10001010_1110_011: DATA = 1'b0;
            15'b10001010_1110_100: DATA = 1'b1;
            15'b10001010_1110_101: DATA = 1'b1;
            15'b10001010_1110_110: DATA = 1'b0;
            15'b10001010_1110_111: DATA = 1'b0;
            // SINE- ROW 0 COL 0 Row 15
            15'b10001010_1111_000: DATA = 1'b0;
            15'b10001010_1111_001: DATA = 1'b0;
            15'b10001010_1111_010: DATA = 1'b0;
            15'b10001010_1111_011: DATA = 1'b0;
            15'b10001010_1111_100: DATA = 1'b0;
            15'b10001010_1111_101: DATA = 1'b1;
            15'b10001010_1111_110: DATA = 1'b0;
            15'b10001010_1111_111: DATA = 1'b0;
            // SINE- ROW 0 COL 1 Row 0
            15'b10001011_0000_000: DATA = 1'b0;
            15'b10001011_0000_001: DATA = 1'b0;
            15'b10001011_0000_010: DATA = 1'b0;
            15'b10001011_0000_011: DATA = 1'b0;
            15'b10001011_0000_100: DATA = 1'b0;
            15'b10001011_0000_101: DATA = 1'b0;
            15'b10001011_0000_110: DATA = 1'b0;
            15'b10001011_0000_111: DATA = 1'b0;
            // SINE- ROW 0 COL 1 Row 1
            15'b10001011_0001_000: DATA = 1'b0;
            15'b10001011_0001_001: DATA = 1'b0;
            15'b10001011_0001_010: DATA = 1'b0;
            15'b10001011_0001_011: DATA = 1'b0;
            15'b10001011_0001_100: DATA = 1'b0;
            15'b10001011_0001_101: DATA = 1'b0;
            15'b10001011_0001_110: DATA = 1'b0;
            15'b10001011_0001_111: DATA = 1'b0;
            // SINE- ROW 0 COL 1 Row 2
            15'b10001011_0010_000: DATA = 1'b0;
            15'b10001011_0010_001: DATA = 1'b0;
            15'b10001011_0010_010: DATA = 1'b0;
            15'b10001011_0010_011: DATA = 1'b0;
            15'b10001011_0010_100: DATA = 1'b0;
            15'b10001011_0010_101: DATA = 1'b0;
            15'b10001011_0010_110: DATA = 1'b0;
            15'b10001011_0010_111: DATA = 1'b0;
            // SINE- ROW 0 COL 1 Row 3
            15'b10001011_0011_000: DATA = 1'b0;
            15'b10001011_0011_001: DATA = 1'b0;
            15'b10001011_0011_010: DATA = 1'b0;
            15'b10001011_0011_011: DATA = 1'b0;
            15'b10001011_0011_100: DATA = 1'b0;
            15'b10001011_0011_101: DATA = 1'b0;
            15'b10001011_0011_110: DATA = 1'b0;
            15'b10001011_0011_111: DATA = 1'b0;
            // SINE- ROW 0 COL 1 Row 4
            15'b10001011_0100_000: DATA = 1'b0;
            15'b10001011_0100_001: DATA = 1'b0;
            15'b10001011_0100_010: DATA = 1'b0;
            15'b10001011_0100_011: DATA = 1'b0;
            15'b10001011_0100_100: DATA = 1'b0;
            15'b10001011_0100_101: DATA = 1'b0;
            15'b10001011_0100_110: DATA = 1'b0;
            15'b10001011_0100_111: DATA = 1'b0;
            // SINE- ROW 0 COL 1 Row 5
            15'b10001011_0101_000: DATA = 1'b0;
            15'b10001011_0101_001: DATA = 1'b0;
            15'b10001011_0101_010: DATA = 1'b0;
            15'b10001011_0101_011: DATA = 1'b0;
            15'b10001011_0101_100: DATA = 1'b0;
            15'b10001011_0101_101: DATA = 1'b0;
            15'b10001011_0101_110: DATA = 1'b0;
            15'b10001011_0101_111: DATA = 1'b0;
            // SINE- ROW 0 COL 1 Row 6
            15'b10001011_0110_000: DATA = 1'b0;
            15'b10001011_0110_001: DATA = 1'b0;
            15'b10001011_0110_010: DATA = 1'b0;
            15'b10001011_0110_011: DATA = 1'b0;
            15'b10001011_0110_100: DATA = 1'b0;
            15'b10001011_0110_101: DATA = 1'b0;
            15'b10001011_0110_110: DATA = 1'b0;
            15'b10001011_0110_111: DATA = 1'b0;
            // SINE- ROW 0 COL 1 Row 7
            15'b10001011_0111_000: DATA = 1'b0;
            15'b10001011_0111_001: DATA = 1'b0;
            15'b10001011_0111_010: DATA = 1'b0;
            15'b10001011_0111_011: DATA = 1'b0;
            15'b10001011_0111_100: DATA = 1'b0;
            15'b10001011_0111_101: DATA = 1'b0;
            15'b10001011_0111_110: DATA = 1'b0;
            15'b10001011_0111_111: DATA = 1'b0;
            // SINE- ROW 0 COL 1 Row 8
            15'b10001011_1000_000: DATA = 1'b0;
            15'b10001011_1000_001: DATA = 1'b0;
            15'b10001011_1000_010: DATA = 1'b0;
            15'b10001011_1000_011: DATA = 1'b0;
            15'b10001011_1000_100: DATA = 1'b0;
            15'b10001011_1000_101: DATA = 1'b0;
            15'b10001011_1000_110: DATA = 1'b0;
            15'b10001011_1000_111: DATA = 1'b0;
            // SINE- ROW 0 COL 1 Row 9
            15'b10001011_1001_000: DATA = 1'b0;
            15'b10001011_1001_001: DATA = 1'b0;
            15'b10001011_1001_010: DATA = 1'b0;
            15'b10001011_1001_011: DATA = 1'b0;
            15'b10001011_1001_100: DATA = 1'b0;
            15'b10001011_1001_101: DATA = 1'b0;
            15'b10001011_1001_110: DATA = 1'b0;
            15'b10001011_1001_111: DATA = 1'b0;
            // SINE- ROW 0 COL 1 Row 10
            15'b10001011_1010_000: DATA = 1'b0;
            15'b10001011_1010_001: DATA = 1'b0;
            15'b10001011_1010_010: DATA = 1'b0;
            15'b10001011_1010_011: DATA = 1'b0;
            15'b10001011_1010_100: DATA = 1'b0;
            15'b10001011_1010_101: DATA = 1'b0;
            15'b10001011_1010_110: DATA = 1'b0;
            15'b10001011_1010_111: DATA = 1'b0;
            // SINE- ROW 0 COL 1 Row 11
            15'b10001011_1011_000: DATA = 1'b0;
            15'b10001011_1011_001: DATA = 1'b0;
            15'b10001011_1011_010: DATA = 1'b0;
            15'b10001011_1011_011: DATA = 1'b0;
            15'b10001011_1011_100: DATA = 1'b0;
            15'b10001011_1011_101: DATA = 1'b0;
            15'b10001011_1011_110: DATA = 1'b0;
            15'b10001011_1011_111: DATA = 1'b0;
            // SINE- ROW 0 COL 1 Row 12
            15'b10001011_1100_000: DATA = 1'b0;
            15'b10001011_1100_001: DATA = 1'b0;
            15'b10001011_1100_010: DATA = 1'b0;
            15'b10001011_1100_011: DATA = 1'b0;
            15'b10001011_1100_100: DATA = 1'b0;
            15'b10001011_1100_101: DATA = 1'b0;
            15'b10001011_1100_110: DATA = 1'b0;
            15'b10001011_1100_111: DATA = 1'b0;
            // SINE- ROW 0 COL 1 Row 13
            15'b10001011_1101_000: DATA = 1'b0;
            15'b10001011_1101_001: DATA = 1'b0;
            15'b10001011_1101_010: DATA = 1'b0;
            15'b10001011_1101_011: DATA = 1'b0;
            15'b10001011_1101_100: DATA = 1'b0;
            15'b10001011_1101_101: DATA = 1'b0;
            15'b10001011_1101_110: DATA = 1'b0;
            15'b10001011_1101_111: DATA = 1'b0;
            // SINE- ROW 0 COL 1 Row 14
            15'b10001011_1110_000: DATA = 1'b0;
            15'b10001011_1110_001: DATA = 1'b0;
            15'b10001011_1110_010: DATA = 1'b0;
            15'b10001011_1110_011: DATA = 1'b0;
            15'b10001011_1110_100: DATA = 1'b0;
            15'b10001011_1110_101: DATA = 1'b0;
            15'b10001011_1110_110: DATA = 1'b0;
            15'b10001011_1110_111: DATA = 1'b0;
            // SINE- ROW 0 COL 1 Row 15
            15'b10001011_1111_000: DATA = 1'b0;
            15'b10001011_1111_001: DATA = 1'b0;
            15'b10001011_1111_010: DATA = 1'b0;
            15'b10001011_1111_011: DATA = 1'b0;
            15'b10001011_1111_100: DATA = 1'b0;
            15'b10001011_1111_101: DATA = 1'b0;
            15'b10001011_1111_110: DATA = 1'b0;
            15'b10001011_1111_111: DATA = 1'b0;
            // SINE- ROW 0 COL 2 Row 0
            15'b10001100_0000_000: DATA = 1'b0;
            15'b10001100_0000_001: DATA = 1'b0;
            15'b10001100_0000_010: DATA = 1'b0;
            15'b10001100_0000_011: DATA = 1'b0;
            15'b10001100_0000_100: DATA = 1'b0;
            15'b10001100_0000_101: DATA = 1'b0;
            15'b10001100_0000_110: DATA = 1'b0;
            15'b10001100_0000_111: DATA = 1'b0;
            // SINE- ROW 0 COL 2 Row 1
            15'b10001100_0001_000: DATA = 1'b0;
            15'b10001100_0001_001: DATA = 1'b0;
            15'b10001100_0001_010: DATA = 1'b0;
            15'b10001100_0001_011: DATA = 1'b0;
            15'b10001100_0001_100: DATA = 1'b0;
            15'b10001100_0001_101: DATA = 1'b0;
            15'b10001100_0001_110: DATA = 1'b0;
            15'b10001100_0001_111: DATA = 1'b0;
            // SINE- ROW 0 COL 2 Row 2
            15'b10001100_0010_000: DATA = 1'b0;
            15'b10001100_0010_001: DATA = 1'b0;
            15'b10001100_0010_010: DATA = 1'b0;
            15'b10001100_0010_011: DATA = 1'b0;
            15'b10001100_0010_100: DATA = 1'b0;
            15'b10001100_0010_101: DATA = 1'b0;
            15'b10001100_0010_110: DATA = 1'b0;
            15'b10001100_0010_111: DATA = 1'b0;
            // SINE- ROW 0 COL 2 Row 3
            15'b10001100_0011_000: DATA = 1'b0;
            15'b10001100_0011_001: DATA = 1'b0;
            15'b10001100_0011_010: DATA = 1'b0;
            15'b10001100_0011_011: DATA = 1'b0;
            15'b10001100_0011_100: DATA = 1'b0;
            15'b10001100_0011_101: DATA = 1'b0;
            15'b10001100_0011_110: DATA = 1'b0;
            15'b10001100_0011_111: DATA = 1'b0;
            // SINE- ROW 0 COL 2 Row 4
            15'b10001100_0100_000: DATA = 1'b0;
            15'b10001100_0100_001: DATA = 1'b0;
            15'b10001100_0100_010: DATA = 1'b0;
            15'b10001100_0100_011: DATA = 1'b0;
            15'b10001100_0100_100: DATA = 1'b0;
            15'b10001100_0100_101: DATA = 1'b0;
            15'b10001100_0100_110: DATA = 1'b0;
            15'b10001100_0100_111: DATA = 1'b0;
            // SINE- ROW 0 COL 2 Row 5
            15'b10001100_0101_000: DATA = 1'b0;
            15'b10001100_0101_001: DATA = 1'b0;
            15'b10001100_0101_010: DATA = 1'b0;
            15'b10001100_0101_011: DATA = 1'b0;
            15'b10001100_0101_100: DATA = 1'b0;
            15'b10001100_0101_101: DATA = 1'b0;
            15'b10001100_0101_110: DATA = 1'b0;
            15'b10001100_0101_111: DATA = 1'b0;
            // SINE- ROW 0 COL 2 Row 6
            15'b10001100_0110_000: DATA = 1'b0;
            15'b10001100_0110_001: DATA = 1'b0;
            15'b10001100_0110_010: DATA = 1'b0;
            15'b10001100_0110_011: DATA = 1'b0;
            15'b10001100_0110_100: DATA = 1'b0;
            15'b10001100_0110_101: DATA = 1'b0;
            15'b10001100_0110_110: DATA = 1'b0;
            15'b10001100_0110_111: DATA = 1'b0;
            // SINE- ROW 0 COL 2 Row 7
            15'b10001100_0111_000: DATA = 1'b0;
            15'b10001100_0111_001: DATA = 1'b0;
            15'b10001100_0111_010: DATA = 1'b0;
            15'b10001100_0111_011: DATA = 1'b0;
            15'b10001100_0111_100: DATA = 1'b0;
            15'b10001100_0111_101: DATA = 1'b0;
            15'b10001100_0111_110: DATA = 1'b0;
            15'b10001100_0111_111: DATA = 1'b0;
            // SINE- ROW 0 COL 2 Row 8
            15'b10001100_1000_000: DATA = 1'b0;
            15'b10001100_1000_001: DATA = 1'b0;
            15'b10001100_1000_010: DATA = 1'b0;
            15'b10001100_1000_011: DATA = 1'b0;
            15'b10001100_1000_100: DATA = 1'b0;
            15'b10001100_1000_101: DATA = 1'b0;
            15'b10001100_1000_110: DATA = 1'b0;
            15'b10001100_1000_111: DATA = 1'b0;
            // SINE- ROW 0 COL 2 Row 9
            15'b10001100_1001_000: DATA = 1'b0;
            15'b10001100_1001_001: DATA = 1'b0;
            15'b10001100_1001_010: DATA = 1'b0;
            15'b10001100_1001_011: DATA = 1'b0;
            15'b10001100_1001_100: DATA = 1'b0;
            15'b10001100_1001_101: DATA = 1'b0;
            15'b10001100_1001_110: DATA = 1'b0;
            15'b10001100_1001_111: DATA = 1'b0;
            // SINE- ROW 0 COL 2 Row 10
            15'b10001100_1010_000: DATA = 1'b0;
            15'b10001100_1010_001: DATA = 1'b0;
            15'b10001100_1010_010: DATA = 1'b0;
            15'b10001100_1010_011: DATA = 1'b0;
            15'b10001100_1010_100: DATA = 1'b0;
            15'b10001100_1010_101: DATA = 1'b0;
            15'b10001100_1010_110: DATA = 1'b0;
            15'b10001100_1010_111: DATA = 1'b0;
            // SINE- ROW 0 COL 2 Row 11
            15'b10001100_1011_000: DATA = 1'b0;
            15'b10001100_1011_001: DATA = 1'b0;
            15'b10001100_1011_010: DATA = 1'b0;
            15'b10001100_1011_011: DATA = 1'b0;
            15'b10001100_1011_100: DATA = 1'b0;
            15'b10001100_1011_101: DATA = 1'b0;
            15'b10001100_1011_110: DATA = 1'b0;
            15'b10001100_1011_111: DATA = 1'b0;
            // SINE- ROW 0 COL 2 Row 12
            15'b10001100_1100_000: DATA = 1'b0;
            15'b10001100_1100_001: DATA = 1'b0;
            15'b10001100_1100_010: DATA = 1'b0;
            15'b10001100_1100_011: DATA = 1'b0;
            15'b10001100_1100_100: DATA = 1'b0;
            15'b10001100_1100_101: DATA = 1'b0;
            15'b10001100_1100_110: DATA = 1'b0;
            15'b10001100_1100_111: DATA = 1'b0;
            // SINE- ROW 0 COL 2 Row 13
            15'b10001100_1101_000: DATA = 1'b0;
            15'b10001100_1101_001: DATA = 1'b0;
            15'b10001100_1101_010: DATA = 1'b0;
            15'b10001100_1101_011: DATA = 1'b0;
            15'b10001100_1101_100: DATA = 1'b0;
            15'b10001100_1101_101: DATA = 1'b0;
            15'b10001100_1101_110: DATA = 1'b0;
            15'b10001100_1101_111: DATA = 1'b0;
            // SINE- ROW 0 COL 2 Row 14
            15'b10001100_1110_000: DATA = 1'b0;
            15'b10001100_1110_001: DATA = 1'b0;
            15'b10001100_1110_010: DATA = 1'b0;
            15'b10001100_1110_011: DATA = 1'b0;
            15'b10001100_1110_100: DATA = 1'b0;
            15'b10001100_1110_101: DATA = 1'b0;
            15'b10001100_1110_110: DATA = 1'b0;
            15'b10001100_1110_111: DATA = 1'b0;
            // SINE- ROW 0 COL 2 Row 15
            15'b10001100_1111_000: DATA = 1'b0;
            15'b10001100_1111_001: DATA = 1'b0;
            15'b10001100_1111_010: DATA = 1'b0;
            15'b10001100_1111_011: DATA = 1'b0;
            15'b10001100_1111_100: DATA = 1'b0;
            15'b10001100_1111_101: DATA = 1'b0;
            15'b10001100_1111_110: DATA = 1'b0;
            15'b10001100_1111_111: DATA = 1'b0;
            // SINE- ROW 0 COL 3 Row 0
            15'b10001101_0000_000: DATA = 1'b0;
            15'b10001101_0000_001: DATA = 1'b0;
            15'b10001101_0000_010: DATA = 1'b0;
            15'b10001101_0000_011: DATA = 1'b0;
            15'b10001101_0000_100: DATA = 1'b0;
            15'b10001101_0000_101: DATA = 1'b0;
            15'b10001101_0000_110: DATA = 1'b0;
            15'b10001101_0000_111: DATA = 1'b0;
            // SINE- ROW 0 COL 3 Row 1
            15'b10001101_0001_000: DATA = 1'b0;
            15'b10001101_0001_001: DATA = 1'b0;
            15'b10001101_0001_010: DATA = 1'b0;
            15'b10001101_0001_011: DATA = 1'b0;
            15'b10001101_0001_100: DATA = 1'b0;
            15'b10001101_0001_101: DATA = 1'b0;
            15'b10001101_0001_110: DATA = 1'b0;
            15'b10001101_0001_111: DATA = 1'b0;
            // SINE- ROW 0 COL 3 Row 2
            15'b10001101_0010_000: DATA = 1'b0;
            15'b10001101_0010_001: DATA = 1'b0;
            15'b10001101_0010_010: DATA = 1'b0;
            15'b10001101_0010_011: DATA = 1'b0;
            15'b10001101_0010_100: DATA = 1'b0;
            15'b10001101_0010_101: DATA = 1'b0;
            15'b10001101_0010_110: DATA = 1'b0;
            15'b10001101_0010_111: DATA = 1'b0;
            // SINE- ROW 0 COL 3 Row 3
            15'b10001101_0011_000: DATA = 1'b0;
            15'b10001101_0011_001: DATA = 1'b0;
            15'b10001101_0011_010: DATA = 1'b0;
            15'b10001101_0011_011: DATA = 1'b0;
            15'b10001101_0011_100: DATA = 1'b0;
            15'b10001101_0011_101: DATA = 1'b0;
            15'b10001101_0011_110: DATA = 1'b0;
            15'b10001101_0011_111: DATA = 1'b0;
            // SINE- ROW 0 COL 3 Row 4
            15'b10001101_0100_000: DATA = 1'b0;
            15'b10001101_0100_001: DATA = 1'b0;
            15'b10001101_0100_010: DATA = 1'b0;
            15'b10001101_0100_011: DATA = 1'b0;
            15'b10001101_0100_100: DATA = 1'b0;
            15'b10001101_0100_101: DATA = 1'b0;
            15'b10001101_0100_110: DATA = 1'b0;
            15'b10001101_0100_111: DATA = 1'b0;
            // SINE- ROW 0 COL 3 Row 5
            15'b10001101_0101_000: DATA = 1'b0;
            15'b10001101_0101_001: DATA = 1'b0;
            15'b10001101_0101_010: DATA = 1'b0;
            15'b10001101_0101_011: DATA = 1'b0;
            15'b10001101_0101_100: DATA = 1'b0;
            15'b10001101_0101_101: DATA = 1'b0;
            15'b10001101_0101_110: DATA = 1'b0;
            15'b10001101_0101_111: DATA = 1'b0;
            // SINE- ROW 0 COL 3 Row 6
            15'b10001101_0110_000: DATA = 1'b0;
            15'b10001101_0110_001: DATA = 1'b0;
            15'b10001101_0110_010: DATA = 1'b0;
            15'b10001101_0110_011: DATA = 1'b0;
            15'b10001101_0110_100: DATA = 1'b0;
            15'b10001101_0110_101: DATA = 1'b0;
            15'b10001101_0110_110: DATA = 1'b0;
            15'b10001101_0110_111: DATA = 1'b0;
            // SINE- ROW 0 COL 3 Row 7
            15'b10001101_0111_000: DATA = 1'b0;
            15'b10001101_0111_001: DATA = 1'b0;
            15'b10001101_0111_010: DATA = 1'b0;
            15'b10001101_0111_011: DATA = 1'b0;
            15'b10001101_0111_100: DATA = 1'b0;
            15'b10001101_0111_101: DATA = 1'b0;
            15'b10001101_0111_110: DATA = 1'b0;
            15'b10001101_0111_111: DATA = 1'b0;
            // SINE- ROW 0 COL 3 Row 8
            15'b10001101_1000_000: DATA = 1'b0;
            15'b10001101_1000_001: DATA = 1'b0;
            15'b10001101_1000_010: DATA = 1'b0;
            15'b10001101_1000_011: DATA = 1'b0;
            15'b10001101_1000_100: DATA = 1'b0;
            15'b10001101_1000_101: DATA = 1'b0;
            15'b10001101_1000_110: DATA = 1'b0;
            15'b10001101_1000_111: DATA = 1'b0;
            // SINE- ROW 0 COL 3 Row 9
            15'b10001101_1001_000: DATA = 1'b0;
            15'b10001101_1001_001: DATA = 1'b0;
            15'b10001101_1001_010: DATA = 1'b0;
            15'b10001101_1001_011: DATA = 1'b0;
            15'b10001101_1001_100: DATA = 1'b0;
            15'b10001101_1001_101: DATA = 1'b0;
            15'b10001101_1001_110: DATA = 1'b0;
            15'b10001101_1001_111: DATA = 1'b0;
            // SINE- ROW 0 COL 3 Row 10
            15'b10001101_1010_000: DATA = 1'b0;
            15'b10001101_1010_001: DATA = 1'b0;
            15'b10001101_1010_010: DATA = 1'b0;
            15'b10001101_1010_011: DATA = 1'b0;
            15'b10001101_1010_100: DATA = 1'b0;
            15'b10001101_1010_101: DATA = 1'b0;
            15'b10001101_1010_110: DATA = 1'b0;
            15'b10001101_1010_111: DATA = 1'b0;
            // SINE- ROW 0 COL 3 Row 11
            15'b10001101_1011_000: DATA = 1'b0;
            15'b10001101_1011_001: DATA = 1'b0;
            15'b10001101_1011_010: DATA = 1'b0;
            15'b10001101_1011_011: DATA = 1'b0;
            15'b10001101_1011_100: DATA = 1'b0;
            15'b10001101_1011_101: DATA = 1'b0;
            15'b10001101_1011_110: DATA = 1'b0;
            15'b10001101_1011_111: DATA = 1'b0;
            // SINE- ROW 0 COL 3 Row 12
            15'b10001101_1100_000: DATA = 1'b0;
            15'b10001101_1100_001: DATA = 1'b0;
            15'b10001101_1100_010: DATA = 1'b0;
            15'b10001101_1100_011: DATA = 1'b0;
            15'b10001101_1100_100: DATA = 1'b0;
            15'b10001101_1100_101: DATA = 1'b0;
            15'b10001101_1100_110: DATA = 1'b0;
            15'b10001101_1100_111: DATA = 1'b0;
            // SINE- ROW 0 COL 3 Row 13
            15'b10001101_1101_000: DATA = 1'b0;
            15'b10001101_1101_001: DATA = 1'b0;
            15'b10001101_1101_010: DATA = 1'b0;
            15'b10001101_1101_011: DATA = 1'b0;
            15'b10001101_1101_100: DATA = 1'b0;
            15'b10001101_1101_101: DATA = 1'b0;
            15'b10001101_1101_110: DATA = 1'b0;
            15'b10001101_1101_111: DATA = 1'b0;
            // SINE- ROW 0 COL 3 Row 14
            15'b10001101_1110_000: DATA = 1'b0;
            15'b10001101_1110_001: DATA = 1'b0;
            15'b10001101_1110_010: DATA = 1'b0;
            15'b10001101_1110_011: DATA = 1'b0;
            15'b10001101_1110_100: DATA = 1'b0;
            15'b10001101_1110_101: DATA = 1'b0;
            15'b10001101_1110_110: DATA = 1'b0;
            15'b10001101_1110_111: DATA = 1'b0;
            // SINE- ROW 0 COL 3 Row 15
            15'b10001101_1111_000: DATA = 1'b0;
            15'b10001101_1111_001: DATA = 1'b0;
            15'b10001101_1111_010: DATA = 1'b0;
            15'b10001101_1111_011: DATA = 1'b0;
            15'b10001101_1111_100: DATA = 1'b0;
            15'b10001101_1111_101: DATA = 1'b0;
            15'b10001101_1111_110: DATA = 1'b0;
            15'b10001101_1111_111: DATA = 1'b0;
            // SINE- ROW 0 COL 4 Row 0
            15'b10001110_0000_000: DATA = 1'b0;
            15'b10001110_0000_001: DATA = 1'b0;
            15'b10001110_0000_010: DATA = 1'b0;
            15'b10001110_0000_011: DATA = 1'b0;
            15'b10001110_0000_100: DATA = 1'b0;
            15'b10001110_0000_101: DATA = 1'b0;
            15'b10001110_0000_110: DATA = 1'b0;
            15'b10001110_0000_111: DATA = 1'b1;
            // SINE- ROW 0 COL 4 Row 1
            15'b10001110_0001_000: DATA = 1'b0;
            15'b10001110_0001_001: DATA = 1'b0;
            15'b10001110_0001_010: DATA = 1'b0;
            15'b10001110_0001_011: DATA = 1'b0;
            15'b10001110_0001_100: DATA = 1'b0;
            15'b10001110_0001_101: DATA = 1'b0;
            15'b10001110_0001_110: DATA = 1'b0;
            15'b10001110_0001_111: DATA = 1'b1;
            // SINE- ROW 0 COL 4 Row 2
            15'b10001110_0010_000: DATA = 1'b0;
            15'b10001110_0010_001: DATA = 1'b0;
            15'b10001110_0010_010: DATA = 1'b0;
            15'b10001110_0010_011: DATA = 1'b0;
            15'b10001110_0010_100: DATA = 1'b0;
            15'b10001110_0010_101: DATA = 1'b0;
            15'b10001110_0010_110: DATA = 1'b0;
            15'b10001110_0010_111: DATA = 1'b1;
            // SINE- ROW 0 COL 4 Row 3
            15'b10001110_0011_000: DATA = 1'b0;
            15'b10001110_0011_001: DATA = 1'b0;
            15'b10001110_0011_010: DATA = 1'b0;
            15'b10001110_0011_011: DATA = 1'b0;
            15'b10001110_0011_100: DATA = 1'b0;
            15'b10001110_0011_101: DATA = 1'b0;
            15'b10001110_0011_110: DATA = 1'b1;
            15'b10001110_0011_111: DATA = 1'b1;
            // SINE- ROW 0 COL 4 Row 4
            15'b10001110_0100_000: DATA = 1'b0;
            15'b10001110_0100_001: DATA = 1'b0;
            15'b10001110_0100_010: DATA = 1'b0;
            15'b10001110_0100_011: DATA = 1'b0;
            15'b10001110_0100_100: DATA = 1'b0;
            15'b10001110_0100_101: DATA = 1'b0;
            15'b10001110_0100_110: DATA = 1'b1;
            15'b10001110_0100_111: DATA = 1'b0;
            // SINE- ROW 0 COL 4 Row 5
            15'b10001110_0101_000: DATA = 1'b0;
            15'b10001110_0101_001: DATA = 1'b0;
            15'b10001110_0101_010: DATA = 1'b0;
            15'b10001110_0101_011: DATA = 1'b0;
            15'b10001110_0101_100: DATA = 1'b0;
            15'b10001110_0101_101: DATA = 1'b0;
            15'b10001110_0101_110: DATA = 1'b1;
            15'b10001110_0101_111: DATA = 1'b0;
            // SINE- ROW 0 COL 4 Row 6
            15'b10001110_0110_000: DATA = 1'b0;
            15'b10001110_0110_001: DATA = 1'b0;
            15'b10001110_0110_010: DATA = 1'b0;
            15'b10001110_0110_011: DATA = 1'b0;
            15'b10001110_0110_100: DATA = 1'b0;
            15'b10001110_0110_101: DATA = 1'b1;
            15'b10001110_0110_110: DATA = 1'b1;
            15'b10001110_0110_111: DATA = 1'b0;
            // SINE- ROW 0 COL 4 Row 7
            15'b10001110_0111_000: DATA = 1'b0;
            15'b10001110_0111_001: DATA = 1'b0;
            15'b10001110_0111_010: DATA = 1'b0;
            15'b10001110_0111_011: DATA = 1'b0;
            15'b10001110_0111_100: DATA = 1'b0;
            15'b10001110_0111_101: DATA = 1'b1;
            15'b10001110_0111_110: DATA = 1'b0;
            15'b10001110_0111_111: DATA = 1'b0;
            // SINE- ROW 0 COL 4 Row 8
            15'b10001110_1000_000: DATA = 1'b0;
            15'b10001110_1000_001: DATA = 1'b0;
            15'b10001110_1000_010: DATA = 1'b0;
            15'b10001110_1000_011: DATA = 1'b0;
            15'b10001110_1000_100: DATA = 1'b0;
            15'b10001110_1000_101: DATA = 1'b1;
            15'b10001110_1000_110: DATA = 1'b0;
            15'b10001110_1000_111: DATA = 1'b0;
            // SINE- ROW 0 COL 4 Row 9
            15'b10001110_1001_000: DATA = 1'b0;
            15'b10001110_1001_001: DATA = 1'b0;
            15'b10001110_1001_010: DATA = 1'b0;
            15'b10001110_1001_011: DATA = 1'b0;
            15'b10001110_1001_100: DATA = 1'b1;
            15'b10001110_1001_101: DATA = 1'b1;
            15'b10001110_1001_110: DATA = 1'b0;
            15'b10001110_1001_111: DATA = 1'b0;
            // SINE- ROW 0 COL 4 Row 10
            15'b10001110_1010_000: DATA = 1'b0;
            15'b10001110_1010_001: DATA = 1'b0;
            15'b10001110_1010_010: DATA = 1'b0;
            15'b10001110_1010_011: DATA = 1'b0;
            15'b10001110_1010_100: DATA = 1'b1;
            15'b10001110_1010_101: DATA = 1'b0;
            15'b10001110_1010_110: DATA = 1'b0;
            15'b10001110_1010_111: DATA = 1'b0;
            // SINE- ROW 0 COL 4 Row 11
            15'b10001110_1011_000: DATA = 1'b0;
            15'b10001110_1011_001: DATA = 1'b0;
            15'b10001110_1011_010: DATA = 1'b0;
            15'b10001110_1011_011: DATA = 1'b0;
            15'b10001110_1011_100: DATA = 1'b1;
            15'b10001110_1011_101: DATA = 1'b0;
            15'b10001110_1011_110: DATA = 1'b0;
            15'b10001110_1011_111: DATA = 1'b0;
            // SINE- ROW 0 COL 4 Row 12
            15'b10001110_1100_000: DATA = 1'b0;
            15'b10001110_1100_001: DATA = 1'b0;
            15'b10001110_1100_010: DATA = 1'b0;
            15'b10001110_1100_011: DATA = 1'b1;
            15'b10001110_1100_100: DATA = 1'b1;
            15'b10001110_1100_101: DATA = 1'b0;
            15'b10001110_1100_110: DATA = 1'b0;
            15'b10001110_1100_111: DATA = 1'b0;
            // SINE- ROW 0 COL 4 Row 13
            15'b10001110_1101_000: DATA = 1'b0;
            15'b10001110_1101_001: DATA = 1'b0;
            15'b10001110_1101_010: DATA = 1'b0;
            15'b10001110_1101_011: DATA = 1'b1;
            15'b10001110_1101_100: DATA = 1'b0;
            15'b10001110_1101_101: DATA = 1'b0;
            15'b10001110_1101_110: DATA = 1'b0;
            15'b10001110_1101_111: DATA = 1'b0;
            // SINE- ROW 0 COL 4 Row 14
            15'b10001110_1110_000: DATA = 1'b0;
            15'b10001110_1110_001: DATA = 1'b0;
            15'b10001110_1110_010: DATA = 1'b1;
            15'b10001110_1110_011: DATA = 1'b1;
            15'b10001110_1110_100: DATA = 1'b0;
            15'b10001110_1110_101: DATA = 1'b0;
            15'b10001110_1110_110: DATA = 1'b0;
            15'b10001110_1110_111: DATA = 1'b0;
            // SINE- ROW 0 COL 4 Row 15
            15'b10001110_1111_000: DATA = 1'b0;
            15'b10001110_1111_001: DATA = 1'b0;
            15'b10001110_1111_010: DATA = 1'b1;
            15'b10001110_1111_011: DATA = 1'b0;
            15'b10001110_1111_100: DATA = 1'b0;
            15'b10001110_1111_101: DATA = 1'b0;
            15'b10001110_1111_110: DATA = 1'b0;
            15'b10001110_1111_111: DATA = 1'b0;
            // SINE- ROW 1 COL 0 Row 0
            15'b10001111_0000_000: DATA = 1'b0;
            15'b10001111_0000_001: DATA = 1'b0;
            15'b10001111_0000_010: DATA = 1'b0;
            15'b10001111_0000_011: DATA = 1'b0;
            15'b10001111_0000_100: DATA = 1'b0;
            15'b10001111_0000_101: DATA = 1'b1;
            15'b10001111_0000_110: DATA = 1'b1;
            15'b10001111_0000_111: DATA = 1'b0;
            // SINE- ROW 1 COL 0 Row 1
            15'b10001111_0001_000: DATA = 1'b0;
            15'b10001111_0001_001: DATA = 1'b0;
            15'b10001111_0001_010: DATA = 1'b0;
            15'b10001111_0001_011: DATA = 1'b0;
            15'b10001111_0001_100: DATA = 1'b0;
            15'b10001111_0001_101: DATA = 1'b0;
            15'b10001111_0001_110: DATA = 1'b1;
            15'b10001111_0001_111: DATA = 1'b0;
            // SINE- ROW 1 COL 0 Row 2
            15'b10001111_0010_000: DATA = 1'b0;
            15'b10001111_0010_001: DATA = 1'b0;
            15'b10001111_0010_010: DATA = 1'b0;
            15'b10001111_0010_011: DATA = 1'b0;
            15'b10001111_0010_100: DATA = 1'b0;
            15'b10001111_0010_101: DATA = 1'b0;
            15'b10001111_0010_110: DATA = 1'b1;
            15'b10001111_0010_111: DATA = 1'b1;
            // SINE- ROW 1 COL 0 Row 3
            15'b10001111_0011_000: DATA = 1'b0;
            15'b10001111_0011_001: DATA = 1'b0;
            15'b10001111_0011_010: DATA = 1'b0;
            15'b10001111_0011_011: DATA = 1'b0;
            15'b10001111_0011_100: DATA = 1'b0;
            15'b10001111_0011_101: DATA = 1'b0;
            15'b10001111_0011_110: DATA = 1'b0;
            15'b10001111_0011_111: DATA = 1'b1;
            // SINE- ROW 1 COL 0 Row 4
            15'b10001111_0100_000: DATA = 1'b0;
            15'b10001111_0100_001: DATA = 1'b0;
            15'b10001111_0100_010: DATA = 1'b0;
            15'b10001111_0100_011: DATA = 1'b0;
            15'b10001111_0100_100: DATA = 1'b0;
            15'b10001111_0100_101: DATA = 1'b0;
            15'b10001111_0100_110: DATA = 1'b0;
            15'b10001111_0100_111: DATA = 1'b1;
            // SINE- ROW 1 COL 0 Row 5
            15'b10001111_0101_000: DATA = 1'b0;
            15'b10001111_0101_001: DATA = 1'b0;
            15'b10001111_0101_010: DATA = 1'b0;
            15'b10001111_0101_011: DATA = 1'b0;
            15'b10001111_0101_100: DATA = 1'b0;
            15'b10001111_0101_101: DATA = 1'b0;
            15'b10001111_0101_110: DATA = 1'b0;
            15'b10001111_0101_111: DATA = 1'b0;
            // SINE- ROW 1 COL 0 Row 6
            15'b10001111_0110_000: DATA = 1'b0;
            15'b10001111_0110_001: DATA = 1'b0;
            15'b10001111_0110_010: DATA = 1'b0;
            15'b10001111_0110_011: DATA = 1'b0;
            15'b10001111_0110_100: DATA = 1'b0;
            15'b10001111_0110_101: DATA = 1'b0;
            15'b10001111_0110_110: DATA = 1'b0;
            15'b10001111_0110_111: DATA = 1'b0;
            // SINE- ROW 1 COL 0 Row 7
            15'b10001111_0111_000: DATA = 1'b0;
            15'b10001111_0111_001: DATA = 1'b0;
            15'b10001111_0111_010: DATA = 1'b0;
            15'b10001111_0111_011: DATA = 1'b0;
            15'b10001111_0111_100: DATA = 1'b0;
            15'b10001111_0111_101: DATA = 1'b0;
            15'b10001111_0111_110: DATA = 1'b0;
            15'b10001111_0111_111: DATA = 1'b0;
            // SINE- ROW 1 COL 0 Row 8
            15'b10001111_1000_000: DATA = 1'b0;
            15'b10001111_1000_001: DATA = 1'b0;
            15'b10001111_1000_010: DATA = 1'b0;
            15'b10001111_1000_011: DATA = 1'b0;
            15'b10001111_1000_100: DATA = 1'b0;
            15'b10001111_1000_101: DATA = 1'b0;
            15'b10001111_1000_110: DATA = 1'b0;
            15'b10001111_1000_111: DATA = 1'b0;
            // SINE- ROW 1 COL 0 Row 9
            15'b10001111_1001_000: DATA = 1'b0;
            15'b10001111_1001_001: DATA = 1'b0;
            15'b10001111_1001_010: DATA = 1'b0;
            15'b10001111_1001_011: DATA = 1'b0;
            15'b10001111_1001_100: DATA = 1'b0;
            15'b10001111_1001_101: DATA = 1'b0;
            15'b10001111_1001_110: DATA = 1'b0;
            15'b10001111_1001_111: DATA = 1'b0;
            // SINE- ROW 1 COL 0 Row 10
            15'b10001111_1010_000: DATA = 1'b0;
            15'b10001111_1010_001: DATA = 1'b0;
            15'b10001111_1010_010: DATA = 1'b0;
            15'b10001111_1010_011: DATA = 1'b0;
            15'b10001111_1010_100: DATA = 1'b0;
            15'b10001111_1010_101: DATA = 1'b0;
            15'b10001111_1010_110: DATA = 1'b0;
            15'b10001111_1010_111: DATA = 1'b0;
            // SINE- ROW 1 COL 0 Row 11
            15'b10001111_1011_000: DATA = 1'b0;
            15'b10001111_1011_001: DATA = 1'b0;
            15'b10001111_1011_010: DATA = 1'b0;
            15'b10001111_1011_011: DATA = 1'b0;
            15'b10001111_1011_100: DATA = 1'b0;
            15'b10001111_1011_101: DATA = 1'b0;
            15'b10001111_1011_110: DATA = 1'b0;
            15'b10001111_1011_111: DATA = 1'b0;
            // SINE- ROW 1 COL 0 Row 12
            15'b10001111_1100_000: DATA = 1'b0;
            15'b10001111_1100_001: DATA = 1'b0;
            15'b10001111_1100_010: DATA = 1'b0;
            15'b10001111_1100_011: DATA = 1'b0;
            15'b10001111_1100_100: DATA = 1'b0;
            15'b10001111_1100_101: DATA = 1'b0;
            15'b10001111_1100_110: DATA = 1'b0;
            15'b10001111_1100_111: DATA = 1'b0;
            // SINE- ROW 1 COL 0 Row 13
            15'b10001111_1101_000: DATA = 1'b0;
            15'b10001111_1101_001: DATA = 1'b0;
            15'b10001111_1101_010: DATA = 1'b0;
            15'b10001111_1101_011: DATA = 1'b0;
            15'b10001111_1101_100: DATA = 1'b0;
            15'b10001111_1101_101: DATA = 1'b0;
            15'b10001111_1101_110: DATA = 1'b0;
            15'b10001111_1101_111: DATA = 1'b0;
            // SINE- ROW 1 COL 0 Row 14
            15'b10001111_1110_000: DATA = 1'b0;
            15'b10001111_1110_001: DATA = 1'b0;
            15'b10001111_1110_010: DATA = 1'b0;
            15'b10001111_1110_011: DATA = 1'b0;
            15'b10001111_1110_100: DATA = 1'b0;
            15'b10001111_1110_101: DATA = 1'b0;
            15'b10001111_1110_110: DATA = 1'b0;
            15'b10001111_1110_111: DATA = 1'b0;
            // SINE- ROW 1 COL 0 Row 15
            15'b10001111_1111_000: DATA = 1'b0;
            15'b10001111_1111_001: DATA = 1'b0;
            15'b10001111_1111_010: DATA = 1'b0;
            15'b10001111_1111_011: DATA = 1'b0;
            15'b10001111_1111_100: DATA = 1'b0;
            15'b10001111_1111_101: DATA = 1'b0;
            15'b10001111_1111_110: DATA = 1'b0;
            15'b10001111_1111_111: DATA = 1'b0;
            // SINE- ROW 1 COL 1 Row 0
            15'b10010000_0000_000: DATA = 1'b0;
            15'b10010000_0000_001: DATA = 1'b0;
            15'b10010000_0000_010: DATA = 1'b0;
            15'b10010000_0000_011: DATA = 1'b0;
            15'b10010000_0000_100: DATA = 1'b0;
            15'b10010000_0000_101: DATA = 1'b0;
            15'b10010000_0000_110: DATA = 1'b0;
            15'b10010000_0000_111: DATA = 1'b0;
            // SINE- ROW 1 COL 1 Row 1
            15'b10010000_0001_000: DATA = 1'b0;
            15'b10010000_0001_001: DATA = 1'b0;
            15'b10010000_0001_010: DATA = 1'b0;
            15'b10010000_0001_011: DATA = 1'b0;
            15'b10010000_0001_100: DATA = 1'b0;
            15'b10010000_0001_101: DATA = 1'b0;
            15'b10010000_0001_110: DATA = 1'b0;
            15'b10010000_0001_111: DATA = 1'b0;
            // SINE- ROW 1 COL 1 Row 2
            15'b10010000_0010_000: DATA = 1'b0;
            15'b10010000_0010_001: DATA = 1'b0;
            15'b10010000_0010_010: DATA = 1'b0;
            15'b10010000_0010_011: DATA = 1'b0;
            15'b10010000_0010_100: DATA = 1'b0;
            15'b10010000_0010_101: DATA = 1'b0;
            15'b10010000_0010_110: DATA = 1'b0;
            15'b10010000_0010_111: DATA = 1'b0;
            // SINE- ROW 1 COL 1 Row 3
            15'b10010000_0011_000: DATA = 1'b0;
            15'b10010000_0011_001: DATA = 1'b0;
            15'b10010000_0011_010: DATA = 1'b0;
            15'b10010000_0011_011: DATA = 1'b0;
            15'b10010000_0011_100: DATA = 1'b0;
            15'b10010000_0011_101: DATA = 1'b0;
            15'b10010000_0011_110: DATA = 1'b0;
            15'b10010000_0011_111: DATA = 1'b0;
            // SINE- ROW 1 COL 1 Row 4
            15'b10010000_0100_000: DATA = 1'b1;
            15'b10010000_0100_001: DATA = 1'b0;
            15'b10010000_0100_010: DATA = 1'b0;
            15'b10010000_0100_011: DATA = 1'b0;
            15'b10010000_0100_100: DATA = 1'b0;
            15'b10010000_0100_101: DATA = 1'b0;
            15'b10010000_0100_110: DATA = 1'b0;
            15'b10010000_0100_111: DATA = 1'b0;
            // SINE- ROW 1 COL 1 Row 5
            15'b10010000_0101_000: DATA = 1'b1;
            15'b10010000_0101_001: DATA = 1'b0;
            15'b10010000_0101_010: DATA = 1'b0;
            15'b10010000_0101_011: DATA = 1'b0;
            15'b10010000_0101_100: DATA = 1'b0;
            15'b10010000_0101_101: DATA = 1'b0;
            15'b10010000_0101_110: DATA = 1'b0;
            15'b10010000_0101_111: DATA = 1'b0;
            // SINE- ROW 1 COL 1 Row 6
            15'b10010000_0110_000: DATA = 1'b1;
            15'b10010000_0110_001: DATA = 1'b1;
            15'b10010000_0110_010: DATA = 1'b0;
            15'b10010000_0110_011: DATA = 1'b0;
            15'b10010000_0110_100: DATA = 1'b0;
            15'b10010000_0110_101: DATA = 1'b0;
            15'b10010000_0110_110: DATA = 1'b0;
            15'b10010000_0110_111: DATA = 1'b0;
            // SINE- ROW 1 COL 1 Row 7
            15'b10010000_0111_000: DATA = 1'b0;
            15'b10010000_0111_001: DATA = 1'b1;
            15'b10010000_0111_010: DATA = 1'b0;
            15'b10010000_0111_011: DATA = 1'b0;
            15'b10010000_0111_100: DATA = 1'b0;
            15'b10010000_0111_101: DATA = 1'b0;
            15'b10010000_0111_110: DATA = 1'b0;
            15'b10010000_0111_111: DATA = 1'b0;
            // SINE- ROW 1 COL 1 Row 8
            15'b10010000_1000_000: DATA = 1'b0;
            15'b10010000_1000_001: DATA = 1'b1;
            15'b10010000_1000_010: DATA = 1'b1;
            15'b10010000_1000_011: DATA = 1'b0;
            15'b10010000_1000_100: DATA = 1'b0;
            15'b10010000_1000_101: DATA = 1'b0;
            15'b10010000_1000_110: DATA = 1'b0;
            15'b10010000_1000_111: DATA = 1'b0;
            // SINE- ROW 1 COL 1 Row 9
            15'b10010000_1001_000: DATA = 1'b0;
            15'b10010000_1001_001: DATA = 1'b0;
            15'b10010000_1001_010: DATA = 1'b1;
            15'b10010000_1001_011: DATA = 1'b1;
            15'b10010000_1001_100: DATA = 1'b0;
            15'b10010000_1001_101: DATA = 1'b0;
            15'b10010000_1001_110: DATA = 1'b0;
            15'b10010000_1001_111: DATA = 1'b0;
            // SINE- ROW 1 COL 1 Row 10
            15'b10010000_1010_000: DATA = 1'b0;
            15'b10010000_1010_001: DATA = 1'b0;
            15'b10010000_1010_010: DATA = 1'b0;
            15'b10010000_1010_011: DATA = 1'b1;
            15'b10010000_1010_100: DATA = 1'b1;
            15'b10010000_1010_101: DATA = 1'b0;
            15'b10010000_1010_110: DATA = 1'b0;
            15'b10010000_1010_111: DATA = 1'b0;
            // SINE- ROW 1 COL 1 Row 11
            15'b10010000_1011_000: DATA = 1'b0;
            15'b10010000_1011_001: DATA = 1'b0;
            15'b10010000_1011_010: DATA = 1'b0;
            15'b10010000_1011_011: DATA = 1'b0;
            15'b10010000_1011_100: DATA = 1'b1;
            15'b10010000_1011_101: DATA = 1'b1;
            15'b10010000_1011_110: DATA = 1'b0;
            15'b10010000_1011_111: DATA = 1'b0;
            // SINE- ROW 1 COL 1 Row 12
            15'b10010000_1100_000: DATA = 1'b0;
            15'b10010000_1100_001: DATA = 1'b0;
            15'b10010000_1100_010: DATA = 1'b0;
            15'b10010000_1100_011: DATA = 1'b0;
            15'b10010000_1100_100: DATA = 1'b0;
            15'b10010000_1100_101: DATA = 1'b1;
            15'b10010000_1100_110: DATA = 1'b1;
            15'b10010000_1100_111: DATA = 1'b0;
            // SINE- ROW 1 COL 1 Row 13
            15'b10010000_1101_000: DATA = 1'b0;
            15'b10010000_1101_001: DATA = 1'b0;
            15'b10010000_1101_010: DATA = 1'b0;
            15'b10010000_1101_011: DATA = 1'b0;
            15'b10010000_1101_100: DATA = 1'b0;
            15'b10010000_1101_101: DATA = 1'b0;
            15'b10010000_1101_110: DATA = 1'b1;
            15'b10010000_1101_111: DATA = 1'b1;
            // SINE- ROW 1 COL 1 Row 14
            15'b10010000_1110_000: DATA = 1'b0;
            15'b10010000_1110_001: DATA = 1'b0;
            15'b10010000_1110_010: DATA = 1'b0;
            15'b10010000_1110_011: DATA = 1'b0;
            15'b10010000_1110_100: DATA = 1'b0;
            15'b10010000_1110_101: DATA = 1'b0;
            15'b10010000_1110_110: DATA = 1'b0;
            15'b10010000_1110_111: DATA = 1'b0;
            // SINE- ROW 1 COL 1 Row 15
            15'b10010000_1111_000: DATA = 1'b0;
            15'b10010000_1111_001: DATA = 1'b0;
            15'b10010000_1111_010: DATA = 1'b0;
            15'b10010000_1111_011: DATA = 1'b0;
            15'b10010000_1111_100: DATA = 1'b0;
            15'b10010000_1111_101: DATA = 1'b0;
            15'b10010000_1111_110: DATA = 1'b0;
            15'b10010000_1111_111: DATA = 1'b0;
            // SINE- ROW 1 COL 2 Row 0
            15'b10010001_0000_000: DATA = 1'b0;
            15'b10010001_0000_001: DATA = 1'b0;
            15'b10010001_0000_010: DATA = 1'b0;
            15'b10010001_0000_011: DATA = 1'b0;
            15'b10010001_0000_100: DATA = 1'b0;
            15'b10010001_0000_101: DATA = 1'b0;
            15'b10010001_0000_110: DATA = 1'b0;
            15'b10010001_0000_111: DATA = 1'b0;
            // SINE- ROW 1 COL 2 Row 1
            15'b10010001_0001_000: DATA = 1'b0;
            15'b10010001_0001_001: DATA = 1'b0;
            15'b10010001_0001_010: DATA = 1'b0;
            15'b10010001_0001_011: DATA = 1'b0;
            15'b10010001_0001_100: DATA = 1'b0;
            15'b10010001_0001_101: DATA = 1'b0;
            15'b10010001_0001_110: DATA = 1'b0;
            15'b10010001_0001_111: DATA = 1'b0;
            // SINE- ROW 1 COL 2 Row 2
            15'b10010001_0010_000: DATA = 1'b0;
            15'b10010001_0010_001: DATA = 1'b0;
            15'b10010001_0010_010: DATA = 1'b0;
            15'b10010001_0010_011: DATA = 1'b0;
            15'b10010001_0010_100: DATA = 1'b0;
            15'b10010001_0010_101: DATA = 1'b0;
            15'b10010001_0010_110: DATA = 1'b0;
            15'b10010001_0010_111: DATA = 1'b0;
            // SINE- ROW 1 COL 2 Row 3
            15'b10010001_0011_000: DATA = 1'b0;
            15'b10010001_0011_001: DATA = 1'b0;
            15'b10010001_0011_010: DATA = 1'b0;
            15'b10010001_0011_011: DATA = 1'b0;
            15'b10010001_0011_100: DATA = 1'b0;
            15'b10010001_0011_101: DATA = 1'b0;
            15'b10010001_0011_110: DATA = 1'b0;
            15'b10010001_0011_111: DATA = 1'b0;
            // SINE- ROW 1 COL 2 Row 4
            15'b10010001_0100_000: DATA = 1'b0;
            15'b10010001_0100_001: DATA = 1'b0;
            15'b10010001_0100_010: DATA = 1'b0;
            15'b10010001_0100_011: DATA = 1'b0;
            15'b10010001_0100_100: DATA = 1'b0;
            15'b10010001_0100_101: DATA = 1'b0;
            15'b10010001_0100_110: DATA = 1'b0;
            15'b10010001_0100_111: DATA = 1'b0;
            // SINE- ROW 1 COL 2 Row 5
            15'b10010001_0101_000: DATA = 1'b0;
            15'b10010001_0101_001: DATA = 1'b0;
            15'b10010001_0101_010: DATA = 1'b0;
            15'b10010001_0101_011: DATA = 1'b0;
            15'b10010001_0101_100: DATA = 1'b0;
            15'b10010001_0101_101: DATA = 1'b0;
            15'b10010001_0101_110: DATA = 1'b0;
            15'b10010001_0101_111: DATA = 1'b0;
            // SINE- ROW 1 COL 2 Row 6
            15'b10010001_0110_000: DATA = 1'b0;
            15'b10010001_0110_001: DATA = 1'b0;
            15'b10010001_0110_010: DATA = 1'b0;
            15'b10010001_0110_011: DATA = 1'b0;
            15'b10010001_0110_100: DATA = 1'b0;
            15'b10010001_0110_101: DATA = 1'b0;
            15'b10010001_0110_110: DATA = 1'b0;
            15'b10010001_0110_111: DATA = 1'b0;
            // SINE- ROW 1 COL 2 Row 7
            15'b10010001_0111_000: DATA = 1'b0;
            15'b10010001_0111_001: DATA = 1'b0;
            15'b10010001_0111_010: DATA = 1'b0;
            15'b10010001_0111_011: DATA = 1'b0;
            15'b10010001_0111_100: DATA = 1'b0;
            15'b10010001_0111_101: DATA = 1'b0;
            15'b10010001_0111_110: DATA = 1'b0;
            15'b10010001_0111_111: DATA = 1'b0;
            // SINE- ROW 1 COL 2 Row 8
            15'b10010001_1000_000: DATA = 1'b0;
            15'b10010001_1000_001: DATA = 1'b0;
            15'b10010001_1000_010: DATA = 1'b0;
            15'b10010001_1000_011: DATA = 1'b0;
            15'b10010001_1000_100: DATA = 1'b0;
            15'b10010001_1000_101: DATA = 1'b0;
            15'b10010001_1000_110: DATA = 1'b0;
            15'b10010001_1000_111: DATA = 1'b0;
            // SINE- ROW 1 COL 2 Row 9
            15'b10010001_1001_000: DATA = 1'b0;
            15'b10010001_1001_001: DATA = 1'b0;
            15'b10010001_1001_010: DATA = 1'b0;
            15'b10010001_1001_011: DATA = 1'b0;
            15'b10010001_1001_100: DATA = 1'b0;
            15'b10010001_1001_101: DATA = 1'b0;
            15'b10010001_1001_110: DATA = 1'b0;
            15'b10010001_1001_111: DATA = 1'b0;
            // SINE- ROW 1 COL 2 Row 10
            15'b10010001_1010_000: DATA = 1'b0;
            15'b10010001_1010_001: DATA = 1'b0;
            15'b10010001_1010_010: DATA = 1'b0;
            15'b10010001_1010_011: DATA = 1'b0;
            15'b10010001_1010_100: DATA = 1'b0;
            15'b10010001_1010_101: DATA = 1'b0;
            15'b10010001_1010_110: DATA = 1'b0;
            15'b10010001_1010_111: DATA = 1'b0;
            // SINE- ROW 1 COL 2 Row 11
            15'b10010001_1011_000: DATA = 1'b0;
            15'b10010001_1011_001: DATA = 1'b0;
            15'b10010001_1011_010: DATA = 1'b0;
            15'b10010001_1011_011: DATA = 1'b0;
            15'b10010001_1011_100: DATA = 1'b0;
            15'b10010001_1011_101: DATA = 1'b0;
            15'b10010001_1011_110: DATA = 1'b0;
            15'b10010001_1011_111: DATA = 1'b0;
            // SINE- ROW 1 COL 2 Row 12
            15'b10010001_1100_000: DATA = 1'b0;
            15'b10010001_1100_001: DATA = 1'b0;
            15'b10010001_1100_010: DATA = 1'b0;
            15'b10010001_1100_011: DATA = 1'b0;
            15'b10010001_1100_100: DATA = 1'b0;
            15'b10010001_1100_101: DATA = 1'b0;
            15'b10010001_1100_110: DATA = 1'b0;
            15'b10010001_1100_111: DATA = 1'b0;
            // SINE- ROW 1 COL 2 Row 13
            15'b10010001_1101_000: DATA = 1'b1;
            15'b10010001_1101_001: DATA = 1'b0;
            15'b10010001_1101_010: DATA = 1'b0;
            15'b10010001_1101_011: DATA = 1'b0;
            15'b10010001_1101_100: DATA = 1'b0;
            15'b10010001_1101_101: DATA = 1'b0;
            15'b10010001_1101_110: DATA = 1'b0;
            15'b10010001_1101_111: DATA = 1'b1;
            // SINE- ROW 1 COL 2 Row 14
            15'b10010001_1110_000: DATA = 1'b1;
            15'b10010001_1110_001: DATA = 1'b1;
            15'b10010001_1110_010: DATA = 1'b1;
            15'b10010001_1110_011: DATA = 1'b0;
            15'b10010001_1110_100: DATA = 1'b0;
            15'b10010001_1110_101: DATA = 1'b1;
            15'b10010001_1110_110: DATA = 1'b1;
            15'b10010001_1110_111: DATA = 1'b1;
            // SINE- ROW 1 COL 2 Row 15
            15'b10010001_1111_000: DATA = 1'b0;
            15'b10010001_1111_001: DATA = 1'b0;
            15'b10010001_1111_010: DATA = 1'b1;
            15'b10010001_1111_011: DATA = 1'b1;
            15'b10010001_1111_100: DATA = 1'b1;
            15'b10010001_1111_101: DATA = 1'b1;
            15'b10010001_1111_110: DATA = 1'b0;
            15'b10010001_1111_111: DATA = 1'b0;
            // SINE- ROW 1 COL 3 Row 0
            15'b10010010_0000_000: DATA = 1'b0;
            15'b10010010_0000_001: DATA = 1'b0;
            15'b10010010_0000_010: DATA = 1'b0;
            15'b10010010_0000_011: DATA = 1'b0;
            15'b10010010_0000_100: DATA = 1'b0;
            15'b10010010_0000_101: DATA = 1'b0;
            15'b10010010_0000_110: DATA = 1'b0;
            15'b10010010_0000_111: DATA = 1'b0;
            // SINE- ROW 1 COL 3 Row 1
            15'b10010010_0001_000: DATA = 1'b0;
            15'b10010010_0001_001: DATA = 1'b0;
            15'b10010010_0001_010: DATA = 1'b0;
            15'b10010010_0001_011: DATA = 1'b0;
            15'b10010010_0001_100: DATA = 1'b0;
            15'b10010010_0001_101: DATA = 1'b0;
            15'b10010010_0001_110: DATA = 1'b0;
            15'b10010010_0001_111: DATA = 1'b0;
            // SINE- ROW 1 COL 3 Row 2
            15'b10010010_0010_000: DATA = 1'b0;
            15'b10010010_0010_001: DATA = 1'b0;
            15'b10010010_0010_010: DATA = 1'b0;
            15'b10010010_0010_011: DATA = 1'b0;
            15'b10010010_0010_100: DATA = 1'b0;
            15'b10010010_0010_101: DATA = 1'b0;
            15'b10010010_0010_110: DATA = 1'b0;
            15'b10010010_0010_111: DATA = 1'b0;
            // SINE- ROW 1 COL 3 Row 3
            15'b10010010_0011_000: DATA = 1'b0;
            15'b10010010_0011_001: DATA = 1'b0;
            15'b10010010_0011_010: DATA = 1'b0;
            15'b10010010_0011_011: DATA = 1'b0;
            15'b10010010_0011_100: DATA = 1'b0;
            15'b10010010_0011_101: DATA = 1'b0;
            15'b10010010_0011_110: DATA = 1'b0;
            15'b10010010_0011_111: DATA = 1'b0;
            // SINE- ROW 1 COL 3 Row 4
            15'b10010010_0100_000: DATA = 1'b0;
            15'b10010010_0100_001: DATA = 1'b0;
            15'b10010010_0100_010: DATA = 1'b0;
            15'b10010010_0100_011: DATA = 1'b0;
            15'b10010010_0100_100: DATA = 1'b0;
            15'b10010010_0100_101: DATA = 1'b0;
            15'b10010010_0100_110: DATA = 1'b0;
            15'b10010010_0100_111: DATA = 1'b1;
            // SINE- ROW 1 COL 3 Row 5
            15'b10010010_0101_000: DATA = 1'b0;
            15'b10010010_0101_001: DATA = 1'b0;
            15'b10010010_0101_010: DATA = 1'b0;
            15'b10010010_0101_011: DATA = 1'b0;
            15'b10010010_0101_100: DATA = 1'b0;
            15'b10010010_0101_101: DATA = 1'b0;
            15'b10010010_0101_110: DATA = 1'b0;
            15'b10010010_0101_111: DATA = 1'b1;
            // SINE- ROW 1 COL 3 Row 6
            15'b10010010_0110_000: DATA = 1'b0;
            15'b10010010_0110_001: DATA = 1'b0;
            15'b10010010_0110_010: DATA = 1'b0;
            15'b10010010_0110_011: DATA = 1'b0;
            15'b10010010_0110_100: DATA = 1'b0;
            15'b10010010_0110_101: DATA = 1'b0;
            15'b10010010_0110_110: DATA = 1'b1;
            15'b10010010_0110_111: DATA = 1'b1;
            // SINE- ROW 1 COL 3 Row 7
            15'b10010010_0111_000: DATA = 1'b0;
            15'b10010010_0111_001: DATA = 1'b0;
            15'b10010010_0111_010: DATA = 1'b0;
            15'b10010010_0111_011: DATA = 1'b0;
            15'b10010010_0111_100: DATA = 1'b0;
            15'b10010010_0111_101: DATA = 1'b0;
            15'b10010010_0111_110: DATA = 1'b1;
            15'b10010010_0111_111: DATA = 1'b0;
            // SINE- ROW 1 COL 3 Row 8
            15'b10010010_1000_000: DATA = 1'b0;
            15'b10010010_1000_001: DATA = 1'b0;
            15'b10010010_1000_010: DATA = 1'b0;
            15'b10010010_1000_011: DATA = 1'b0;
            15'b10010010_1000_100: DATA = 1'b0;
            15'b10010010_1000_101: DATA = 1'b1;
            15'b10010010_1000_110: DATA = 1'b1;
            15'b10010010_1000_111: DATA = 1'b0;
            // SINE- ROW 1 COL 3 Row 9
            15'b10010010_1001_000: DATA = 1'b0;
            15'b10010010_1001_001: DATA = 1'b0;
            15'b10010010_1001_010: DATA = 1'b0;
            15'b10010010_1001_011: DATA = 1'b0;
            15'b10010010_1001_100: DATA = 1'b1;
            15'b10010010_1001_101: DATA = 1'b1;
            15'b10010010_1001_110: DATA = 1'b0;
            15'b10010010_1001_111: DATA = 1'b0;
            // SINE- ROW 1 COL 3 Row 10
            15'b10010010_1010_000: DATA = 1'b0;
            15'b10010010_1010_001: DATA = 1'b0;
            15'b10010010_1010_010: DATA = 1'b0;
            15'b10010010_1010_011: DATA = 1'b1;
            15'b10010010_1010_100: DATA = 1'b1;
            15'b10010010_1010_101: DATA = 1'b0;
            15'b10010010_1010_110: DATA = 1'b0;
            15'b10010010_1010_111: DATA = 1'b0;
            // SINE- ROW 1 COL 3 Row 11
            15'b10010010_1011_000: DATA = 1'b0;
            15'b10010010_1011_001: DATA = 1'b0;
            15'b10010010_1011_010: DATA = 1'b1;
            15'b10010010_1011_011: DATA = 1'b1;
            15'b10010010_1011_100: DATA = 1'b0;
            15'b10010010_1011_101: DATA = 1'b0;
            15'b10010010_1011_110: DATA = 1'b0;
            15'b10010010_1011_111: DATA = 1'b0;
            // SINE- ROW 1 COL 3 Row 12
            15'b10010010_1100_000: DATA = 1'b0;
            15'b10010010_1100_001: DATA = 1'b1;
            15'b10010010_1100_010: DATA = 1'b1;
            15'b10010010_1100_011: DATA = 1'b0;
            15'b10010010_1100_100: DATA = 1'b0;
            15'b10010010_1100_101: DATA = 1'b0;
            15'b10010010_1100_110: DATA = 1'b0;
            15'b10010010_1100_111: DATA = 1'b0;
            // SINE- ROW 1 COL 3 Row 13
            15'b10010010_1101_000: DATA = 1'b1;
            15'b10010010_1101_001: DATA = 1'b1;
            15'b10010010_1101_010: DATA = 1'b0;
            15'b10010010_1101_011: DATA = 1'b0;
            15'b10010010_1101_100: DATA = 1'b0;
            15'b10010010_1101_101: DATA = 1'b0;
            15'b10010010_1101_110: DATA = 1'b0;
            15'b10010010_1101_111: DATA = 1'b0;
            // SINE- ROW 1 COL 3 Row 14
            15'b10010010_1110_000: DATA = 1'b0;
            15'b10010010_1110_001: DATA = 1'b0;
            15'b10010010_1110_010: DATA = 1'b0;
            15'b10010010_1110_011: DATA = 1'b0;
            15'b10010010_1110_100: DATA = 1'b0;
            15'b10010010_1110_101: DATA = 1'b0;
            15'b10010010_1110_110: DATA = 1'b0;
            15'b10010010_1110_111: DATA = 1'b0;
            // SINE- ROW 1 COL 3 Row 15
            15'b10010010_1111_000: DATA = 1'b0;
            15'b10010010_1111_001: DATA = 1'b0;
            15'b10010010_1111_010: DATA = 1'b0;
            15'b10010010_1111_011: DATA = 1'b0;
            15'b10010010_1111_100: DATA = 1'b0;
            15'b10010010_1111_101: DATA = 1'b0;
            15'b10010010_1111_110: DATA = 1'b0;
            15'b10010010_1111_111: DATA = 1'b0;
            // SINE- ROW 1 COL 4 Row 0
            15'b10010011_0000_000: DATA = 1'b0;
            15'b10010011_0000_001: DATA = 1'b1;
            15'b10010011_0000_010: DATA = 1'b1;
            15'b10010011_0000_011: DATA = 1'b0;
            15'b10010011_0000_100: DATA = 1'b0;
            15'b10010011_0000_101: DATA = 1'b0;
            15'b10010011_0000_110: DATA = 1'b0;
            15'b10010011_0000_111: DATA = 1'b0;
            // SINE- ROW 1 COL 4 Row 1
            15'b10010011_0001_000: DATA = 1'b0;
            15'b10010011_0001_001: DATA = 1'b1;
            15'b10010011_0001_010: DATA = 1'b0;
            15'b10010011_0001_011: DATA = 1'b0;
            15'b10010011_0001_100: DATA = 1'b0;
            15'b10010011_0001_101: DATA = 1'b0;
            15'b10010011_0001_110: DATA = 1'b0;
            15'b10010011_0001_111: DATA = 1'b0;
            // SINE- ROW 1 COL 4 Row 2
            15'b10010011_0010_000: DATA = 1'b1;
            15'b10010011_0010_001: DATA = 1'b1;
            15'b10010011_0010_010: DATA = 1'b0;
            15'b10010011_0010_011: DATA = 1'b0;
            15'b10010011_0010_100: DATA = 1'b0;
            15'b10010011_0010_101: DATA = 1'b0;
            15'b10010011_0010_110: DATA = 1'b0;
            15'b10010011_0010_111: DATA = 1'b0;
            // SINE- ROW 1 COL 4 Row 3
            15'b10010011_0011_000: DATA = 1'b1;
            15'b10010011_0011_001: DATA = 1'b0;
            15'b10010011_0011_010: DATA = 1'b0;
            15'b10010011_0011_011: DATA = 1'b0;
            15'b10010011_0011_100: DATA = 1'b0;
            15'b10010011_0011_101: DATA = 1'b0;
            15'b10010011_0011_110: DATA = 1'b0;
            15'b10010011_0011_111: DATA = 1'b0;
            // SINE- ROW 1 COL 4 Row 4
            15'b10010011_0100_000: DATA = 1'b1;
            15'b10010011_0100_001: DATA = 1'b0;
            15'b10010011_0100_010: DATA = 1'b0;
            15'b10010011_0100_011: DATA = 1'b0;
            15'b10010011_0100_100: DATA = 1'b0;
            15'b10010011_0100_101: DATA = 1'b0;
            15'b10010011_0100_110: DATA = 1'b0;
            15'b10010011_0100_111: DATA = 1'b0;
            // SINE- ROW 1 COL 4 Row 5
            15'b10010011_0101_000: DATA = 1'b0;
            15'b10010011_0101_001: DATA = 1'b0;
            15'b10010011_0101_010: DATA = 1'b0;
            15'b10010011_0101_011: DATA = 1'b0;
            15'b10010011_0101_100: DATA = 1'b0;
            15'b10010011_0101_101: DATA = 1'b0;
            15'b10010011_0101_110: DATA = 1'b0;
            15'b10010011_0101_111: DATA = 1'b0;
            // SINE- ROW 1 COL 4 Row 6
            15'b10010011_0110_000: DATA = 1'b0;
            15'b10010011_0110_001: DATA = 1'b0;
            15'b10010011_0110_010: DATA = 1'b0;
            15'b10010011_0110_011: DATA = 1'b0;
            15'b10010011_0110_100: DATA = 1'b0;
            15'b10010011_0110_101: DATA = 1'b0;
            15'b10010011_0110_110: DATA = 1'b0;
            15'b10010011_0110_111: DATA = 1'b0;
            // SINE- ROW 1 COL 4 Row 7
            15'b10010011_0111_000: DATA = 1'b0;
            15'b10010011_0111_001: DATA = 1'b0;
            15'b10010011_0111_010: DATA = 1'b0;
            15'b10010011_0111_011: DATA = 1'b0;
            15'b10010011_0111_100: DATA = 1'b0;
            15'b10010011_0111_101: DATA = 1'b0;
            15'b10010011_0111_110: DATA = 1'b0;
            15'b10010011_0111_111: DATA = 1'b0;
            // SINE- ROW 1 COL 4 Row 8
            15'b10010011_1000_000: DATA = 1'b0;
            15'b10010011_1000_001: DATA = 1'b0;
            15'b10010011_1000_010: DATA = 1'b0;
            15'b10010011_1000_011: DATA = 1'b0;
            15'b10010011_1000_100: DATA = 1'b0;
            15'b10010011_1000_101: DATA = 1'b0;
            15'b10010011_1000_110: DATA = 1'b0;
            15'b10010011_1000_111: DATA = 1'b0;
            // SINE- ROW 1 COL 4 Row 9
            15'b10010011_1001_000: DATA = 1'b0;
            15'b10010011_1001_001: DATA = 1'b0;
            15'b10010011_1001_010: DATA = 1'b0;
            15'b10010011_1001_011: DATA = 1'b0;
            15'b10010011_1001_100: DATA = 1'b0;
            15'b10010011_1001_101: DATA = 1'b0;
            15'b10010011_1001_110: DATA = 1'b0;
            15'b10010011_1001_111: DATA = 1'b0;
            // SINE- ROW 1 COL 4 Row 10
            15'b10010011_1010_000: DATA = 1'b0;
            15'b10010011_1010_001: DATA = 1'b0;
            15'b10010011_1010_010: DATA = 1'b0;
            15'b10010011_1010_011: DATA = 1'b0;
            15'b10010011_1010_100: DATA = 1'b0;
            15'b10010011_1010_101: DATA = 1'b0;
            15'b10010011_1010_110: DATA = 1'b0;
            15'b10010011_1010_111: DATA = 1'b0;
            // SINE- ROW 1 COL 4 Row 11
            15'b10010011_1011_000: DATA = 1'b0;
            15'b10010011_1011_001: DATA = 1'b0;
            15'b10010011_1011_010: DATA = 1'b0;
            15'b10010011_1011_011: DATA = 1'b0;
            15'b10010011_1011_100: DATA = 1'b0;
            15'b10010011_1011_101: DATA = 1'b0;
            15'b10010011_1011_110: DATA = 1'b0;
            15'b10010011_1011_111: DATA = 1'b0;
            // SINE- ROW 1 COL 4 Row 12
            15'b10010011_1100_000: DATA = 1'b0;
            15'b10010011_1100_001: DATA = 1'b0;
            15'b10010011_1100_010: DATA = 1'b0;
            15'b10010011_1100_011: DATA = 1'b0;
            15'b10010011_1100_100: DATA = 1'b0;
            15'b10010011_1100_101: DATA = 1'b0;
            15'b10010011_1100_110: DATA = 1'b0;
            15'b10010011_1100_111: DATA = 1'b0;
            // SINE- ROW 1 COL 4 Row 13
            15'b10010011_1101_000: DATA = 1'b0;
            15'b10010011_1101_001: DATA = 1'b0;
            15'b10010011_1101_010: DATA = 1'b0;
            15'b10010011_1101_011: DATA = 1'b0;
            15'b10010011_1101_100: DATA = 1'b0;
            15'b10010011_1101_101: DATA = 1'b0;
            15'b10010011_1101_110: DATA = 1'b0;
            15'b10010011_1101_111: DATA = 1'b0;
            // SINE- ROW 1 COL 4 Row 14
            15'b10010011_1110_000: DATA = 1'b0;
            15'b10010011_1110_001: DATA = 1'b0;
            15'b10010011_1110_010: DATA = 1'b0;
            15'b10010011_1110_011: DATA = 1'b0;
            15'b10010011_1110_100: DATA = 1'b0;
            15'b10010011_1110_101: DATA = 1'b0;
            15'b10010011_1110_110: DATA = 1'b0;
            15'b10010011_1110_111: DATA = 1'b0;
            // SINE- ROW 1 COL 4 Row 15
            15'b10010011_1111_000: DATA = 1'b0;
            15'b10010011_1111_001: DATA = 1'b0;
            15'b10010011_1111_010: DATA = 1'b0;
            15'b10010011_1111_011: DATA = 1'b0;
            15'b10010011_1111_100: DATA = 1'b0;
            15'b10010011_1111_101: DATA = 1'b0;
            15'b10010011_1111_110: DATA = 1'b0;
            15'b10010011_1111_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 0 Row 0
            15'b10010100_0000_000: DATA = 1'b1;
            15'b10010100_0000_001: DATA = 1'b1;
            15'b10010100_0000_010: DATA = 1'b1;
            15'b10010100_0000_011: DATA = 1'b1;
            15'b10010100_0000_100: DATA = 1'b1;
            15'b10010100_0000_101: DATA = 1'b1;
            15'b10010100_0000_110: DATA = 1'b1;
            15'b10010100_0000_111: DATA = 1'b1;
            // SQUARE+ ROW 0 COL 0 Row 1
            15'b10010100_0001_000: DATA = 1'b1;
            15'b10010100_0001_001: DATA = 1'b0;
            15'b10010100_0001_010: DATA = 1'b0;
            15'b10010100_0001_011: DATA = 1'b0;
            15'b10010100_0001_100: DATA = 1'b0;
            15'b10010100_0001_101: DATA = 1'b0;
            15'b10010100_0001_110: DATA = 1'b0;
            15'b10010100_0001_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 0 Row 2
            15'b10010100_0010_000: DATA = 1'b1;
            15'b10010100_0010_001: DATA = 1'b0;
            15'b10010100_0010_010: DATA = 1'b0;
            15'b10010100_0010_011: DATA = 1'b0;
            15'b10010100_0010_100: DATA = 1'b0;
            15'b10010100_0010_101: DATA = 1'b0;
            15'b10010100_0010_110: DATA = 1'b0;
            15'b10010100_0010_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 0 Row 3
            15'b10010100_0011_000: DATA = 1'b1;
            15'b10010100_0011_001: DATA = 1'b0;
            15'b10010100_0011_010: DATA = 1'b0;
            15'b10010100_0011_011: DATA = 1'b0;
            15'b10010100_0011_100: DATA = 1'b0;
            15'b10010100_0011_101: DATA = 1'b0;
            15'b10010100_0011_110: DATA = 1'b0;
            15'b10010100_0011_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 0 Row 4
            15'b10010100_0100_000: DATA = 1'b1;
            15'b10010100_0100_001: DATA = 1'b0;
            15'b10010100_0100_010: DATA = 1'b0;
            15'b10010100_0100_011: DATA = 1'b0;
            15'b10010100_0100_100: DATA = 1'b0;
            15'b10010100_0100_101: DATA = 1'b0;
            15'b10010100_0100_110: DATA = 1'b0;
            15'b10010100_0100_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 0 Row 5
            15'b10010100_0101_000: DATA = 1'b1;
            15'b10010100_0101_001: DATA = 1'b0;
            15'b10010100_0101_010: DATA = 1'b0;
            15'b10010100_0101_011: DATA = 1'b0;
            15'b10010100_0101_100: DATA = 1'b0;
            15'b10010100_0101_101: DATA = 1'b0;
            15'b10010100_0101_110: DATA = 1'b0;
            15'b10010100_0101_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 0 Row 6
            15'b10010100_0110_000: DATA = 1'b1;
            15'b10010100_0110_001: DATA = 1'b0;
            15'b10010100_0110_010: DATA = 1'b0;
            15'b10010100_0110_011: DATA = 1'b0;
            15'b10010100_0110_100: DATA = 1'b0;
            15'b10010100_0110_101: DATA = 1'b0;
            15'b10010100_0110_110: DATA = 1'b0;
            15'b10010100_0110_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 0 Row 7
            15'b10010100_0111_000: DATA = 1'b1;
            15'b10010100_0111_001: DATA = 1'b0;
            15'b10010100_0111_010: DATA = 1'b0;
            15'b10010100_0111_011: DATA = 1'b0;
            15'b10010100_0111_100: DATA = 1'b0;
            15'b10010100_0111_101: DATA = 1'b0;
            15'b10010100_0111_110: DATA = 1'b0;
            15'b10010100_0111_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 0 Row 8
            15'b10010100_1000_000: DATA = 1'b1;
            15'b10010100_1000_001: DATA = 1'b0;
            15'b10010100_1000_010: DATA = 1'b0;
            15'b10010100_1000_011: DATA = 1'b0;
            15'b10010100_1000_100: DATA = 1'b0;
            15'b10010100_1000_101: DATA = 1'b0;
            15'b10010100_1000_110: DATA = 1'b0;
            15'b10010100_1000_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 0 Row 9
            15'b10010100_1001_000: DATA = 1'b1;
            15'b10010100_1001_001: DATA = 1'b0;
            15'b10010100_1001_010: DATA = 1'b0;
            15'b10010100_1001_011: DATA = 1'b0;
            15'b10010100_1001_100: DATA = 1'b0;
            15'b10010100_1001_101: DATA = 1'b0;
            15'b10010100_1001_110: DATA = 1'b0;
            15'b10010100_1001_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 0 Row 10
            15'b10010100_1010_000: DATA = 1'b1;
            15'b10010100_1010_001: DATA = 1'b0;
            15'b10010100_1010_010: DATA = 1'b0;
            15'b10010100_1010_011: DATA = 1'b0;
            15'b10010100_1010_100: DATA = 1'b0;
            15'b10010100_1010_101: DATA = 1'b0;
            15'b10010100_1010_110: DATA = 1'b0;
            15'b10010100_1010_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 0 Row 11
            15'b10010100_1011_000: DATA = 1'b1;
            15'b10010100_1011_001: DATA = 1'b0;
            15'b10010100_1011_010: DATA = 1'b0;
            15'b10010100_1011_011: DATA = 1'b0;
            15'b10010100_1011_100: DATA = 1'b0;
            15'b10010100_1011_101: DATA = 1'b0;
            15'b10010100_1011_110: DATA = 1'b0;
            15'b10010100_1011_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 0 Row 12
            15'b10010100_1100_000: DATA = 1'b1;
            15'b10010100_1100_001: DATA = 1'b0;
            15'b10010100_1100_010: DATA = 1'b0;
            15'b10010100_1100_011: DATA = 1'b0;
            15'b10010100_1100_100: DATA = 1'b0;
            15'b10010100_1100_101: DATA = 1'b0;
            15'b10010100_1100_110: DATA = 1'b0;
            15'b10010100_1100_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 0 Row 13
            15'b10010100_1101_000: DATA = 1'b1;
            15'b10010100_1101_001: DATA = 1'b0;
            15'b10010100_1101_010: DATA = 1'b0;
            15'b10010100_1101_011: DATA = 1'b0;
            15'b10010100_1101_100: DATA = 1'b0;
            15'b10010100_1101_101: DATA = 1'b0;
            15'b10010100_1101_110: DATA = 1'b0;
            15'b10010100_1101_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 0 Row 14
            15'b10010100_1110_000: DATA = 1'b1;
            15'b10010100_1110_001: DATA = 1'b0;
            15'b10010100_1110_010: DATA = 1'b0;
            15'b10010100_1110_011: DATA = 1'b0;
            15'b10010100_1110_100: DATA = 1'b0;
            15'b10010100_1110_101: DATA = 1'b0;
            15'b10010100_1110_110: DATA = 1'b0;
            15'b10010100_1110_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 0 Row 15
            15'b10010100_1111_000: DATA = 1'b1;
            15'b10010100_1111_001: DATA = 1'b0;
            15'b10010100_1111_010: DATA = 1'b0;
            15'b10010100_1111_011: DATA = 1'b0;
            15'b10010100_1111_100: DATA = 1'b0;
            15'b10010100_1111_101: DATA = 1'b0;
            15'b10010100_1111_110: DATA = 1'b0;
            15'b10010100_1111_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 1 Row 0
            15'b10010101_0000_000: DATA = 1'b1;
            15'b10010101_0000_001: DATA = 1'b1;
            15'b10010101_0000_010: DATA = 1'b1;
            15'b10010101_0000_011: DATA = 1'b1;
            15'b10010101_0000_100: DATA = 1'b1;
            15'b10010101_0000_101: DATA = 1'b1;
            15'b10010101_0000_110: DATA = 1'b1;
            15'b10010101_0000_111: DATA = 1'b1;
            // SQUARE+ ROW 0 COL 1 Row 1
            15'b10010101_0001_000: DATA = 1'b0;
            15'b10010101_0001_001: DATA = 1'b0;
            15'b10010101_0001_010: DATA = 1'b0;
            15'b10010101_0001_011: DATA = 1'b0;
            15'b10010101_0001_100: DATA = 1'b0;
            15'b10010101_0001_101: DATA = 1'b0;
            15'b10010101_0001_110: DATA = 1'b0;
            15'b10010101_0001_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 1 Row 2
            15'b10010101_0010_000: DATA = 1'b0;
            15'b10010101_0010_001: DATA = 1'b0;
            15'b10010101_0010_010: DATA = 1'b0;
            15'b10010101_0010_011: DATA = 1'b0;
            15'b10010101_0010_100: DATA = 1'b0;
            15'b10010101_0010_101: DATA = 1'b0;
            15'b10010101_0010_110: DATA = 1'b0;
            15'b10010101_0010_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 1 Row 3
            15'b10010101_0011_000: DATA = 1'b0;
            15'b10010101_0011_001: DATA = 1'b0;
            15'b10010101_0011_010: DATA = 1'b0;
            15'b10010101_0011_011: DATA = 1'b0;
            15'b10010101_0011_100: DATA = 1'b0;
            15'b10010101_0011_101: DATA = 1'b0;
            15'b10010101_0011_110: DATA = 1'b0;
            15'b10010101_0011_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 1 Row 4
            15'b10010101_0100_000: DATA = 1'b0;
            15'b10010101_0100_001: DATA = 1'b0;
            15'b10010101_0100_010: DATA = 1'b0;
            15'b10010101_0100_011: DATA = 1'b0;
            15'b10010101_0100_100: DATA = 1'b0;
            15'b10010101_0100_101: DATA = 1'b0;
            15'b10010101_0100_110: DATA = 1'b0;
            15'b10010101_0100_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 1 Row 5
            15'b10010101_0101_000: DATA = 1'b0;
            15'b10010101_0101_001: DATA = 1'b0;
            15'b10010101_0101_010: DATA = 1'b0;
            15'b10010101_0101_011: DATA = 1'b0;
            15'b10010101_0101_100: DATA = 1'b0;
            15'b10010101_0101_101: DATA = 1'b0;
            15'b10010101_0101_110: DATA = 1'b0;
            15'b10010101_0101_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 1 Row 6
            15'b10010101_0110_000: DATA = 1'b0;
            15'b10010101_0110_001: DATA = 1'b0;
            15'b10010101_0110_010: DATA = 1'b0;
            15'b10010101_0110_011: DATA = 1'b0;
            15'b10010101_0110_100: DATA = 1'b0;
            15'b10010101_0110_101: DATA = 1'b0;
            15'b10010101_0110_110: DATA = 1'b0;
            15'b10010101_0110_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 1 Row 7
            15'b10010101_0111_000: DATA = 1'b0;
            15'b10010101_0111_001: DATA = 1'b0;
            15'b10010101_0111_010: DATA = 1'b0;
            15'b10010101_0111_011: DATA = 1'b0;
            15'b10010101_0111_100: DATA = 1'b0;
            15'b10010101_0111_101: DATA = 1'b0;
            15'b10010101_0111_110: DATA = 1'b0;
            15'b10010101_0111_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 1 Row 8
            15'b10010101_1000_000: DATA = 1'b0;
            15'b10010101_1000_001: DATA = 1'b0;
            15'b10010101_1000_010: DATA = 1'b0;
            15'b10010101_1000_011: DATA = 1'b0;
            15'b10010101_1000_100: DATA = 1'b0;
            15'b10010101_1000_101: DATA = 1'b0;
            15'b10010101_1000_110: DATA = 1'b0;
            15'b10010101_1000_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 1 Row 9
            15'b10010101_1001_000: DATA = 1'b0;
            15'b10010101_1001_001: DATA = 1'b0;
            15'b10010101_1001_010: DATA = 1'b0;
            15'b10010101_1001_011: DATA = 1'b0;
            15'b10010101_1001_100: DATA = 1'b0;
            15'b10010101_1001_101: DATA = 1'b0;
            15'b10010101_1001_110: DATA = 1'b0;
            15'b10010101_1001_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 1 Row 10
            15'b10010101_1010_000: DATA = 1'b0;
            15'b10010101_1010_001: DATA = 1'b0;
            15'b10010101_1010_010: DATA = 1'b0;
            15'b10010101_1010_011: DATA = 1'b0;
            15'b10010101_1010_100: DATA = 1'b0;
            15'b10010101_1010_101: DATA = 1'b0;
            15'b10010101_1010_110: DATA = 1'b0;
            15'b10010101_1010_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 1 Row 11
            15'b10010101_1011_000: DATA = 1'b0;
            15'b10010101_1011_001: DATA = 1'b0;
            15'b10010101_1011_010: DATA = 1'b0;
            15'b10010101_1011_011: DATA = 1'b0;
            15'b10010101_1011_100: DATA = 1'b0;
            15'b10010101_1011_101: DATA = 1'b0;
            15'b10010101_1011_110: DATA = 1'b0;
            15'b10010101_1011_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 1 Row 12
            15'b10010101_1100_000: DATA = 1'b0;
            15'b10010101_1100_001: DATA = 1'b0;
            15'b10010101_1100_010: DATA = 1'b0;
            15'b10010101_1100_011: DATA = 1'b0;
            15'b10010101_1100_100: DATA = 1'b0;
            15'b10010101_1100_101: DATA = 1'b0;
            15'b10010101_1100_110: DATA = 1'b0;
            15'b10010101_1100_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 1 Row 13
            15'b10010101_1101_000: DATA = 1'b0;
            15'b10010101_1101_001: DATA = 1'b0;
            15'b10010101_1101_010: DATA = 1'b0;
            15'b10010101_1101_011: DATA = 1'b0;
            15'b10010101_1101_100: DATA = 1'b0;
            15'b10010101_1101_101: DATA = 1'b0;
            15'b10010101_1101_110: DATA = 1'b0;
            15'b10010101_1101_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 1 Row 14
            15'b10010101_1110_000: DATA = 1'b0;
            15'b10010101_1110_001: DATA = 1'b0;
            15'b10010101_1110_010: DATA = 1'b0;
            15'b10010101_1110_011: DATA = 1'b0;
            15'b10010101_1110_100: DATA = 1'b0;
            15'b10010101_1110_101: DATA = 1'b0;
            15'b10010101_1110_110: DATA = 1'b0;
            15'b10010101_1110_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 1 Row 15
            15'b10010101_1111_000: DATA = 1'b0;
            15'b10010101_1111_001: DATA = 1'b0;
            15'b10010101_1111_010: DATA = 1'b0;
            15'b10010101_1111_011: DATA = 1'b0;
            15'b10010101_1111_100: DATA = 1'b0;
            15'b10010101_1111_101: DATA = 1'b0;
            15'b10010101_1111_110: DATA = 1'b0;
            15'b10010101_1111_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 2 Row 0
            15'b10010110_0000_000: DATA = 1'b1;
            15'b10010110_0000_001: DATA = 1'b1;
            15'b10010110_0000_010: DATA = 1'b1;
            15'b10010110_0000_011: DATA = 1'b1;
            15'b10010110_0000_100: DATA = 1'b1;
            15'b10010110_0000_101: DATA = 1'b1;
            15'b10010110_0000_110: DATA = 1'b1;
            15'b10010110_0000_111: DATA = 1'b1;
            // SQUARE+ ROW 0 COL 2 Row 1
            15'b10010110_0001_000: DATA = 1'b0;
            15'b10010110_0001_001: DATA = 1'b0;
            15'b10010110_0001_010: DATA = 1'b0;
            15'b10010110_0001_011: DATA = 1'b0;
            15'b10010110_0001_100: DATA = 1'b0;
            15'b10010110_0001_101: DATA = 1'b0;
            15'b10010110_0001_110: DATA = 1'b0;
            15'b10010110_0001_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 2 Row 2
            15'b10010110_0010_000: DATA = 1'b0;
            15'b10010110_0010_001: DATA = 1'b0;
            15'b10010110_0010_010: DATA = 1'b0;
            15'b10010110_0010_011: DATA = 1'b0;
            15'b10010110_0010_100: DATA = 1'b0;
            15'b10010110_0010_101: DATA = 1'b0;
            15'b10010110_0010_110: DATA = 1'b0;
            15'b10010110_0010_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 2 Row 3
            15'b10010110_0011_000: DATA = 1'b0;
            15'b10010110_0011_001: DATA = 1'b0;
            15'b10010110_0011_010: DATA = 1'b0;
            15'b10010110_0011_011: DATA = 1'b0;
            15'b10010110_0011_100: DATA = 1'b0;
            15'b10010110_0011_101: DATA = 1'b0;
            15'b10010110_0011_110: DATA = 1'b0;
            15'b10010110_0011_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 2 Row 4
            15'b10010110_0100_000: DATA = 1'b0;
            15'b10010110_0100_001: DATA = 1'b0;
            15'b10010110_0100_010: DATA = 1'b0;
            15'b10010110_0100_011: DATA = 1'b0;
            15'b10010110_0100_100: DATA = 1'b0;
            15'b10010110_0100_101: DATA = 1'b0;
            15'b10010110_0100_110: DATA = 1'b0;
            15'b10010110_0100_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 2 Row 5
            15'b10010110_0101_000: DATA = 1'b0;
            15'b10010110_0101_001: DATA = 1'b0;
            15'b10010110_0101_010: DATA = 1'b0;
            15'b10010110_0101_011: DATA = 1'b0;
            15'b10010110_0101_100: DATA = 1'b0;
            15'b10010110_0101_101: DATA = 1'b0;
            15'b10010110_0101_110: DATA = 1'b0;
            15'b10010110_0101_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 2 Row 6
            15'b10010110_0110_000: DATA = 1'b0;
            15'b10010110_0110_001: DATA = 1'b0;
            15'b10010110_0110_010: DATA = 1'b0;
            15'b10010110_0110_011: DATA = 1'b0;
            15'b10010110_0110_100: DATA = 1'b0;
            15'b10010110_0110_101: DATA = 1'b0;
            15'b10010110_0110_110: DATA = 1'b0;
            15'b10010110_0110_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 2 Row 7
            15'b10010110_0111_000: DATA = 1'b0;
            15'b10010110_0111_001: DATA = 1'b0;
            15'b10010110_0111_010: DATA = 1'b0;
            15'b10010110_0111_011: DATA = 1'b0;
            15'b10010110_0111_100: DATA = 1'b0;
            15'b10010110_0111_101: DATA = 1'b0;
            15'b10010110_0111_110: DATA = 1'b0;
            15'b10010110_0111_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 2 Row 8
            15'b10010110_1000_000: DATA = 1'b0;
            15'b10010110_1000_001: DATA = 1'b0;
            15'b10010110_1000_010: DATA = 1'b0;
            15'b10010110_1000_011: DATA = 1'b0;
            15'b10010110_1000_100: DATA = 1'b0;
            15'b10010110_1000_101: DATA = 1'b0;
            15'b10010110_1000_110: DATA = 1'b0;
            15'b10010110_1000_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 2 Row 9
            15'b10010110_1001_000: DATA = 1'b0;
            15'b10010110_1001_001: DATA = 1'b0;
            15'b10010110_1001_010: DATA = 1'b0;
            15'b10010110_1001_011: DATA = 1'b0;
            15'b10010110_1001_100: DATA = 1'b0;
            15'b10010110_1001_101: DATA = 1'b0;
            15'b10010110_1001_110: DATA = 1'b0;
            15'b10010110_1001_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 2 Row 10
            15'b10010110_1010_000: DATA = 1'b0;
            15'b10010110_1010_001: DATA = 1'b0;
            15'b10010110_1010_010: DATA = 1'b0;
            15'b10010110_1010_011: DATA = 1'b0;
            15'b10010110_1010_100: DATA = 1'b0;
            15'b10010110_1010_101: DATA = 1'b0;
            15'b10010110_1010_110: DATA = 1'b0;
            15'b10010110_1010_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 2 Row 11
            15'b10010110_1011_000: DATA = 1'b0;
            15'b10010110_1011_001: DATA = 1'b0;
            15'b10010110_1011_010: DATA = 1'b0;
            15'b10010110_1011_011: DATA = 1'b0;
            15'b10010110_1011_100: DATA = 1'b0;
            15'b10010110_1011_101: DATA = 1'b0;
            15'b10010110_1011_110: DATA = 1'b0;
            15'b10010110_1011_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 2 Row 12
            15'b10010110_1100_000: DATA = 1'b0;
            15'b10010110_1100_001: DATA = 1'b0;
            15'b10010110_1100_010: DATA = 1'b0;
            15'b10010110_1100_011: DATA = 1'b0;
            15'b10010110_1100_100: DATA = 1'b0;
            15'b10010110_1100_101: DATA = 1'b0;
            15'b10010110_1100_110: DATA = 1'b0;
            15'b10010110_1100_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 2 Row 13
            15'b10010110_1101_000: DATA = 1'b0;
            15'b10010110_1101_001: DATA = 1'b0;
            15'b10010110_1101_010: DATA = 1'b0;
            15'b10010110_1101_011: DATA = 1'b0;
            15'b10010110_1101_100: DATA = 1'b0;
            15'b10010110_1101_101: DATA = 1'b0;
            15'b10010110_1101_110: DATA = 1'b0;
            15'b10010110_1101_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 2 Row 14
            15'b10010110_1110_000: DATA = 1'b0;
            15'b10010110_1110_001: DATA = 1'b0;
            15'b10010110_1110_010: DATA = 1'b0;
            15'b10010110_1110_011: DATA = 1'b0;
            15'b10010110_1110_100: DATA = 1'b0;
            15'b10010110_1110_101: DATA = 1'b0;
            15'b10010110_1110_110: DATA = 1'b0;
            15'b10010110_1110_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 2 Row 15
            15'b10010110_1111_000: DATA = 1'b0;
            15'b10010110_1111_001: DATA = 1'b0;
            15'b10010110_1111_010: DATA = 1'b0;
            15'b10010110_1111_011: DATA = 1'b0;
            15'b10010110_1111_100: DATA = 1'b0;
            15'b10010110_1111_101: DATA = 1'b0;
            15'b10010110_1111_110: DATA = 1'b0;
            15'b10010110_1111_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 3 Row 0
            15'b10010111_0000_000: DATA = 1'b1;
            15'b10010111_0000_001: DATA = 1'b1;
            15'b10010111_0000_010: DATA = 1'b1;
            15'b10010111_0000_011: DATA = 1'b1;
            15'b10010111_0000_100: DATA = 1'b1;
            15'b10010111_0000_101: DATA = 1'b1;
            15'b10010111_0000_110: DATA = 1'b1;
            15'b10010111_0000_111: DATA = 1'b1;
            // SQUARE+ ROW 0 COL 3 Row 1
            15'b10010111_0001_000: DATA = 1'b0;
            15'b10010111_0001_001: DATA = 1'b0;
            15'b10010111_0001_010: DATA = 1'b0;
            15'b10010111_0001_011: DATA = 1'b0;
            15'b10010111_0001_100: DATA = 1'b0;
            15'b10010111_0001_101: DATA = 1'b0;
            15'b10010111_0001_110: DATA = 1'b0;
            15'b10010111_0001_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 3 Row 2
            15'b10010111_0010_000: DATA = 1'b0;
            15'b10010111_0010_001: DATA = 1'b0;
            15'b10010111_0010_010: DATA = 1'b0;
            15'b10010111_0010_011: DATA = 1'b0;
            15'b10010111_0010_100: DATA = 1'b0;
            15'b10010111_0010_101: DATA = 1'b0;
            15'b10010111_0010_110: DATA = 1'b0;
            15'b10010111_0010_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 3 Row 3
            15'b10010111_0011_000: DATA = 1'b0;
            15'b10010111_0011_001: DATA = 1'b0;
            15'b10010111_0011_010: DATA = 1'b0;
            15'b10010111_0011_011: DATA = 1'b0;
            15'b10010111_0011_100: DATA = 1'b0;
            15'b10010111_0011_101: DATA = 1'b0;
            15'b10010111_0011_110: DATA = 1'b0;
            15'b10010111_0011_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 3 Row 4
            15'b10010111_0100_000: DATA = 1'b0;
            15'b10010111_0100_001: DATA = 1'b0;
            15'b10010111_0100_010: DATA = 1'b0;
            15'b10010111_0100_011: DATA = 1'b0;
            15'b10010111_0100_100: DATA = 1'b0;
            15'b10010111_0100_101: DATA = 1'b0;
            15'b10010111_0100_110: DATA = 1'b0;
            15'b10010111_0100_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 3 Row 5
            15'b10010111_0101_000: DATA = 1'b0;
            15'b10010111_0101_001: DATA = 1'b0;
            15'b10010111_0101_010: DATA = 1'b0;
            15'b10010111_0101_011: DATA = 1'b0;
            15'b10010111_0101_100: DATA = 1'b0;
            15'b10010111_0101_101: DATA = 1'b0;
            15'b10010111_0101_110: DATA = 1'b0;
            15'b10010111_0101_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 3 Row 6
            15'b10010111_0110_000: DATA = 1'b0;
            15'b10010111_0110_001: DATA = 1'b0;
            15'b10010111_0110_010: DATA = 1'b0;
            15'b10010111_0110_011: DATA = 1'b0;
            15'b10010111_0110_100: DATA = 1'b0;
            15'b10010111_0110_101: DATA = 1'b0;
            15'b10010111_0110_110: DATA = 1'b0;
            15'b10010111_0110_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 3 Row 7
            15'b10010111_0111_000: DATA = 1'b0;
            15'b10010111_0111_001: DATA = 1'b0;
            15'b10010111_0111_010: DATA = 1'b0;
            15'b10010111_0111_011: DATA = 1'b0;
            15'b10010111_0111_100: DATA = 1'b0;
            15'b10010111_0111_101: DATA = 1'b0;
            15'b10010111_0111_110: DATA = 1'b0;
            15'b10010111_0111_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 3 Row 8
            15'b10010111_1000_000: DATA = 1'b0;
            15'b10010111_1000_001: DATA = 1'b0;
            15'b10010111_1000_010: DATA = 1'b0;
            15'b10010111_1000_011: DATA = 1'b0;
            15'b10010111_1000_100: DATA = 1'b0;
            15'b10010111_1000_101: DATA = 1'b0;
            15'b10010111_1000_110: DATA = 1'b0;
            15'b10010111_1000_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 3 Row 9
            15'b10010111_1001_000: DATA = 1'b0;
            15'b10010111_1001_001: DATA = 1'b0;
            15'b10010111_1001_010: DATA = 1'b0;
            15'b10010111_1001_011: DATA = 1'b0;
            15'b10010111_1001_100: DATA = 1'b0;
            15'b10010111_1001_101: DATA = 1'b0;
            15'b10010111_1001_110: DATA = 1'b0;
            15'b10010111_1001_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 3 Row 10
            15'b10010111_1010_000: DATA = 1'b0;
            15'b10010111_1010_001: DATA = 1'b0;
            15'b10010111_1010_010: DATA = 1'b0;
            15'b10010111_1010_011: DATA = 1'b0;
            15'b10010111_1010_100: DATA = 1'b0;
            15'b10010111_1010_101: DATA = 1'b0;
            15'b10010111_1010_110: DATA = 1'b0;
            15'b10010111_1010_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 3 Row 11
            15'b10010111_1011_000: DATA = 1'b0;
            15'b10010111_1011_001: DATA = 1'b0;
            15'b10010111_1011_010: DATA = 1'b0;
            15'b10010111_1011_011: DATA = 1'b0;
            15'b10010111_1011_100: DATA = 1'b0;
            15'b10010111_1011_101: DATA = 1'b0;
            15'b10010111_1011_110: DATA = 1'b0;
            15'b10010111_1011_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 3 Row 12
            15'b10010111_1100_000: DATA = 1'b0;
            15'b10010111_1100_001: DATA = 1'b0;
            15'b10010111_1100_010: DATA = 1'b0;
            15'b10010111_1100_011: DATA = 1'b0;
            15'b10010111_1100_100: DATA = 1'b0;
            15'b10010111_1100_101: DATA = 1'b0;
            15'b10010111_1100_110: DATA = 1'b0;
            15'b10010111_1100_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 3 Row 13
            15'b10010111_1101_000: DATA = 1'b0;
            15'b10010111_1101_001: DATA = 1'b0;
            15'b10010111_1101_010: DATA = 1'b0;
            15'b10010111_1101_011: DATA = 1'b0;
            15'b10010111_1101_100: DATA = 1'b0;
            15'b10010111_1101_101: DATA = 1'b0;
            15'b10010111_1101_110: DATA = 1'b0;
            15'b10010111_1101_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 3 Row 14
            15'b10010111_1110_000: DATA = 1'b0;
            15'b10010111_1110_001: DATA = 1'b0;
            15'b10010111_1110_010: DATA = 1'b0;
            15'b10010111_1110_011: DATA = 1'b0;
            15'b10010111_1110_100: DATA = 1'b0;
            15'b10010111_1110_101: DATA = 1'b0;
            15'b10010111_1110_110: DATA = 1'b0;
            15'b10010111_1110_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 3 Row 15
            15'b10010111_1111_000: DATA = 1'b0;
            15'b10010111_1111_001: DATA = 1'b0;
            15'b10010111_1111_010: DATA = 1'b0;
            15'b10010111_1111_011: DATA = 1'b0;
            15'b10010111_1111_100: DATA = 1'b0;
            15'b10010111_1111_101: DATA = 1'b0;
            15'b10010111_1111_110: DATA = 1'b0;
            15'b10010111_1111_111: DATA = 1'b0;
            // SQUARE+ ROW 0 COL 4 Row 0
            15'b10011000_0000_000: DATA = 1'b1;
            15'b10011000_0000_001: DATA = 1'b1;
            15'b10011000_0000_010: DATA = 1'b1;
            15'b10011000_0000_011: DATA = 1'b1;
            15'b10011000_0000_100: DATA = 1'b1;
            15'b10011000_0000_101: DATA = 1'b1;
            15'b10011000_0000_110: DATA = 1'b1;
            15'b10011000_0000_111: DATA = 1'b1;
            // SQUARE+ ROW 0 COL 4 Row 1
            15'b10011000_0001_000: DATA = 1'b0;
            15'b10011000_0001_001: DATA = 1'b0;
            15'b10011000_0001_010: DATA = 1'b0;
            15'b10011000_0001_011: DATA = 1'b0;
            15'b10011000_0001_100: DATA = 1'b0;
            15'b10011000_0001_101: DATA = 1'b0;
            15'b10011000_0001_110: DATA = 1'b0;
            15'b10011000_0001_111: DATA = 1'b1;
            // SQUARE+ ROW 0 COL 4 Row 2
            15'b10011000_0010_000: DATA = 1'b0;
            15'b10011000_0010_001: DATA = 1'b0;
            15'b10011000_0010_010: DATA = 1'b0;
            15'b10011000_0010_011: DATA = 1'b0;
            15'b10011000_0010_100: DATA = 1'b0;
            15'b10011000_0010_101: DATA = 1'b0;
            15'b10011000_0010_110: DATA = 1'b0;
            15'b10011000_0010_111: DATA = 1'b1;
            // SQUARE+ ROW 0 COL 4 Row 3
            15'b10011000_0011_000: DATA = 1'b0;
            15'b10011000_0011_001: DATA = 1'b0;
            15'b10011000_0011_010: DATA = 1'b0;
            15'b10011000_0011_011: DATA = 1'b0;
            15'b10011000_0011_100: DATA = 1'b0;
            15'b10011000_0011_101: DATA = 1'b0;
            15'b10011000_0011_110: DATA = 1'b0;
            15'b10011000_0011_111: DATA = 1'b1;
            // SQUARE+ ROW 0 COL 4 Row 4
            15'b10011000_0100_000: DATA = 1'b0;
            15'b10011000_0100_001: DATA = 1'b0;
            15'b10011000_0100_010: DATA = 1'b0;
            15'b10011000_0100_011: DATA = 1'b0;
            15'b10011000_0100_100: DATA = 1'b0;
            15'b10011000_0100_101: DATA = 1'b0;
            15'b10011000_0100_110: DATA = 1'b0;
            15'b10011000_0100_111: DATA = 1'b1;
            // SQUARE+ ROW 0 COL 4 Row 5
            15'b10011000_0101_000: DATA = 1'b0;
            15'b10011000_0101_001: DATA = 1'b0;
            15'b10011000_0101_010: DATA = 1'b0;
            15'b10011000_0101_011: DATA = 1'b0;
            15'b10011000_0101_100: DATA = 1'b0;
            15'b10011000_0101_101: DATA = 1'b0;
            15'b10011000_0101_110: DATA = 1'b0;
            15'b10011000_0101_111: DATA = 1'b1;
            // SQUARE+ ROW 0 COL 4 Row 6
            15'b10011000_0110_000: DATA = 1'b0;
            15'b10011000_0110_001: DATA = 1'b0;
            15'b10011000_0110_010: DATA = 1'b0;
            15'b10011000_0110_011: DATA = 1'b0;
            15'b10011000_0110_100: DATA = 1'b0;
            15'b10011000_0110_101: DATA = 1'b0;
            15'b10011000_0110_110: DATA = 1'b0;
            15'b10011000_0110_111: DATA = 1'b1;
            // SQUARE+ ROW 0 COL 4 Row 7
            15'b10011000_0111_000: DATA = 1'b0;
            15'b10011000_0111_001: DATA = 1'b0;
            15'b10011000_0111_010: DATA = 1'b0;
            15'b10011000_0111_011: DATA = 1'b0;
            15'b10011000_0111_100: DATA = 1'b0;
            15'b10011000_0111_101: DATA = 1'b0;
            15'b10011000_0111_110: DATA = 1'b0;
            15'b10011000_0111_111: DATA = 1'b1;
            // SQUARE+ ROW 0 COL 4 Row 8
            15'b10011000_1000_000: DATA = 1'b0;
            15'b10011000_1000_001: DATA = 1'b0;
            15'b10011000_1000_010: DATA = 1'b0;
            15'b10011000_1000_011: DATA = 1'b0;
            15'b10011000_1000_100: DATA = 1'b0;
            15'b10011000_1000_101: DATA = 1'b0;
            15'b10011000_1000_110: DATA = 1'b0;
            15'b10011000_1000_111: DATA = 1'b1;
            // SQUARE+ ROW 0 COL 4 Row 9
            15'b10011000_1001_000: DATA = 1'b0;
            15'b10011000_1001_001: DATA = 1'b0;
            15'b10011000_1001_010: DATA = 1'b0;
            15'b10011000_1001_011: DATA = 1'b0;
            15'b10011000_1001_100: DATA = 1'b0;
            15'b10011000_1001_101: DATA = 1'b0;
            15'b10011000_1001_110: DATA = 1'b0;
            15'b10011000_1001_111: DATA = 1'b1;
            // SQUARE+ ROW 0 COL 4 Row 10
            15'b10011000_1010_000: DATA = 1'b0;
            15'b10011000_1010_001: DATA = 1'b0;
            15'b10011000_1010_010: DATA = 1'b0;
            15'b10011000_1010_011: DATA = 1'b0;
            15'b10011000_1010_100: DATA = 1'b0;
            15'b10011000_1010_101: DATA = 1'b0;
            15'b10011000_1010_110: DATA = 1'b0;
            15'b10011000_1010_111: DATA = 1'b1;
            // SQUARE+ ROW 0 COL 4 Row 11
            15'b10011000_1011_000: DATA = 1'b0;
            15'b10011000_1011_001: DATA = 1'b0;
            15'b10011000_1011_010: DATA = 1'b0;
            15'b10011000_1011_011: DATA = 1'b0;
            15'b10011000_1011_100: DATA = 1'b0;
            15'b10011000_1011_101: DATA = 1'b0;
            15'b10011000_1011_110: DATA = 1'b0;
            15'b10011000_1011_111: DATA = 1'b1;
            // SQUARE+ ROW 0 COL 4 Row 12
            15'b10011000_1100_000: DATA = 1'b0;
            15'b10011000_1100_001: DATA = 1'b0;
            15'b10011000_1100_010: DATA = 1'b0;
            15'b10011000_1100_011: DATA = 1'b0;
            15'b10011000_1100_100: DATA = 1'b0;
            15'b10011000_1100_101: DATA = 1'b0;
            15'b10011000_1100_110: DATA = 1'b0;
            15'b10011000_1100_111: DATA = 1'b1;
            // SQUARE+ ROW 0 COL 4 Row 13
            15'b10011000_1101_000: DATA = 1'b0;
            15'b10011000_1101_001: DATA = 1'b0;
            15'b10011000_1101_010: DATA = 1'b0;
            15'b10011000_1101_011: DATA = 1'b0;
            15'b10011000_1101_100: DATA = 1'b0;
            15'b10011000_1101_101: DATA = 1'b0;
            15'b10011000_1101_110: DATA = 1'b0;
            15'b10011000_1101_111: DATA = 1'b1;
            // SQUARE+ ROW 0 COL 4 Row 14
            15'b10011000_1110_000: DATA = 1'b0;
            15'b10011000_1110_001: DATA = 1'b0;
            15'b10011000_1110_010: DATA = 1'b0;
            15'b10011000_1110_011: DATA = 1'b0;
            15'b10011000_1110_100: DATA = 1'b0;
            15'b10011000_1110_101: DATA = 1'b0;
            15'b10011000_1110_110: DATA = 1'b0;
            15'b10011000_1110_111: DATA = 1'b1;
            // SQUARE+ ROW 0 COL 4 Row 15
            15'b10011000_1111_000: DATA = 1'b0;
            15'b10011000_1111_001: DATA = 1'b0;
            15'b10011000_1111_010: DATA = 1'b0;
            15'b10011000_1111_011: DATA = 1'b0;
            15'b10011000_1111_100: DATA = 1'b0;
            15'b10011000_1111_101: DATA = 1'b0;
            15'b10011000_1111_110: DATA = 1'b0;
            15'b10011000_1111_111: DATA = 1'b1;
            // SQUARE+ ROW 1 COL 0 Row 0
            15'b10011001_0000_000: DATA = 1'b1;
            15'b10011001_0000_001: DATA = 1'b0;
            15'b10011001_0000_010: DATA = 1'b0;
            15'b10011001_0000_011: DATA = 1'b0;
            15'b10011001_0000_100: DATA = 1'b0;
            15'b10011001_0000_101: DATA = 1'b0;
            15'b10011001_0000_110: DATA = 1'b0;
            15'b10011001_0000_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 0 Row 1
            15'b10011001_0001_000: DATA = 1'b1;
            15'b10011001_0001_001: DATA = 1'b0;
            15'b10011001_0001_010: DATA = 1'b0;
            15'b10011001_0001_011: DATA = 1'b0;
            15'b10011001_0001_100: DATA = 1'b0;
            15'b10011001_0001_101: DATA = 1'b0;
            15'b10011001_0001_110: DATA = 1'b0;
            15'b10011001_0001_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 0 Row 2
            15'b10011001_0010_000: DATA = 1'b1;
            15'b10011001_0010_001: DATA = 1'b0;
            15'b10011001_0010_010: DATA = 1'b0;
            15'b10011001_0010_011: DATA = 1'b0;
            15'b10011001_0010_100: DATA = 1'b0;
            15'b10011001_0010_101: DATA = 1'b0;
            15'b10011001_0010_110: DATA = 1'b0;
            15'b10011001_0010_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 0 Row 3
            15'b10011001_0011_000: DATA = 1'b1;
            15'b10011001_0011_001: DATA = 1'b0;
            15'b10011001_0011_010: DATA = 1'b0;
            15'b10011001_0011_011: DATA = 1'b0;
            15'b10011001_0011_100: DATA = 1'b0;
            15'b10011001_0011_101: DATA = 1'b0;
            15'b10011001_0011_110: DATA = 1'b0;
            15'b10011001_0011_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 0 Row 4
            15'b10011001_0100_000: DATA = 1'b1;
            15'b10011001_0100_001: DATA = 1'b0;
            15'b10011001_0100_010: DATA = 1'b0;
            15'b10011001_0100_011: DATA = 1'b0;
            15'b10011001_0100_100: DATA = 1'b0;
            15'b10011001_0100_101: DATA = 1'b0;
            15'b10011001_0100_110: DATA = 1'b0;
            15'b10011001_0100_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 0 Row 5
            15'b10011001_0101_000: DATA = 1'b1;
            15'b10011001_0101_001: DATA = 1'b0;
            15'b10011001_0101_010: DATA = 1'b0;
            15'b10011001_0101_011: DATA = 1'b0;
            15'b10011001_0101_100: DATA = 1'b0;
            15'b10011001_0101_101: DATA = 1'b0;
            15'b10011001_0101_110: DATA = 1'b0;
            15'b10011001_0101_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 0 Row 6
            15'b10011001_0110_000: DATA = 1'b1;
            15'b10011001_0110_001: DATA = 1'b0;
            15'b10011001_0110_010: DATA = 1'b0;
            15'b10011001_0110_011: DATA = 1'b0;
            15'b10011001_0110_100: DATA = 1'b0;
            15'b10011001_0110_101: DATA = 1'b0;
            15'b10011001_0110_110: DATA = 1'b0;
            15'b10011001_0110_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 0 Row 7
            15'b10011001_0111_000: DATA = 1'b1;
            15'b10011001_0111_001: DATA = 1'b0;
            15'b10011001_0111_010: DATA = 1'b0;
            15'b10011001_0111_011: DATA = 1'b0;
            15'b10011001_0111_100: DATA = 1'b0;
            15'b10011001_0111_101: DATA = 1'b0;
            15'b10011001_0111_110: DATA = 1'b0;
            15'b10011001_0111_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 0 Row 8
            15'b10011001_1000_000: DATA = 1'b1;
            15'b10011001_1000_001: DATA = 1'b0;
            15'b10011001_1000_010: DATA = 1'b0;
            15'b10011001_1000_011: DATA = 1'b0;
            15'b10011001_1000_100: DATA = 1'b0;
            15'b10011001_1000_101: DATA = 1'b0;
            15'b10011001_1000_110: DATA = 1'b0;
            15'b10011001_1000_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 0 Row 9
            15'b10011001_1001_000: DATA = 1'b1;
            15'b10011001_1001_001: DATA = 1'b0;
            15'b10011001_1001_010: DATA = 1'b0;
            15'b10011001_1001_011: DATA = 1'b0;
            15'b10011001_1001_100: DATA = 1'b0;
            15'b10011001_1001_101: DATA = 1'b0;
            15'b10011001_1001_110: DATA = 1'b0;
            15'b10011001_1001_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 0 Row 10
            15'b10011001_1010_000: DATA = 1'b1;
            15'b10011001_1010_001: DATA = 1'b0;
            15'b10011001_1010_010: DATA = 1'b0;
            15'b10011001_1010_011: DATA = 1'b0;
            15'b10011001_1010_100: DATA = 1'b0;
            15'b10011001_1010_101: DATA = 1'b0;
            15'b10011001_1010_110: DATA = 1'b0;
            15'b10011001_1010_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 0 Row 11
            15'b10011001_1011_000: DATA = 1'b1;
            15'b10011001_1011_001: DATA = 1'b0;
            15'b10011001_1011_010: DATA = 1'b0;
            15'b10011001_1011_011: DATA = 1'b0;
            15'b10011001_1011_100: DATA = 1'b0;
            15'b10011001_1011_101: DATA = 1'b0;
            15'b10011001_1011_110: DATA = 1'b0;
            15'b10011001_1011_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 0 Row 12
            15'b10011001_1100_000: DATA = 1'b1;
            15'b10011001_1100_001: DATA = 1'b0;
            15'b10011001_1100_010: DATA = 1'b0;
            15'b10011001_1100_011: DATA = 1'b0;
            15'b10011001_1100_100: DATA = 1'b0;
            15'b10011001_1100_101: DATA = 1'b0;
            15'b10011001_1100_110: DATA = 1'b0;
            15'b10011001_1100_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 0 Row 13
            15'b10011001_1101_000: DATA = 1'b1;
            15'b10011001_1101_001: DATA = 1'b0;
            15'b10011001_1101_010: DATA = 1'b0;
            15'b10011001_1101_011: DATA = 1'b0;
            15'b10011001_1101_100: DATA = 1'b0;
            15'b10011001_1101_101: DATA = 1'b0;
            15'b10011001_1101_110: DATA = 1'b0;
            15'b10011001_1101_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 0 Row 14
            15'b10011001_1110_000: DATA = 1'b1;
            15'b10011001_1110_001: DATA = 1'b0;
            15'b10011001_1110_010: DATA = 1'b0;
            15'b10011001_1110_011: DATA = 1'b0;
            15'b10011001_1110_100: DATA = 1'b0;
            15'b10011001_1110_101: DATA = 1'b0;
            15'b10011001_1110_110: DATA = 1'b0;
            15'b10011001_1110_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 0 Row 15
            15'b10011001_1111_000: DATA = 1'b1;
            15'b10011001_1111_001: DATA = 1'b0;
            15'b10011001_1111_010: DATA = 1'b0;
            15'b10011001_1111_011: DATA = 1'b0;
            15'b10011001_1111_100: DATA = 1'b0;
            15'b10011001_1111_101: DATA = 1'b0;
            15'b10011001_1111_110: DATA = 1'b0;
            15'b10011001_1111_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 1 Row 0
            15'b10011010_0000_000: DATA = 1'b0;
            15'b10011010_0000_001: DATA = 1'b0;
            15'b10011010_0000_010: DATA = 1'b0;
            15'b10011010_0000_011: DATA = 1'b0;
            15'b10011010_0000_100: DATA = 1'b0;
            15'b10011010_0000_101: DATA = 1'b0;
            15'b10011010_0000_110: DATA = 1'b0;
            15'b10011010_0000_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 1 Row 1
            15'b10011010_0001_000: DATA = 1'b0;
            15'b10011010_0001_001: DATA = 1'b0;
            15'b10011010_0001_010: DATA = 1'b0;
            15'b10011010_0001_011: DATA = 1'b0;
            15'b10011010_0001_100: DATA = 1'b0;
            15'b10011010_0001_101: DATA = 1'b0;
            15'b10011010_0001_110: DATA = 1'b0;
            15'b10011010_0001_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 1 Row 2
            15'b10011010_0010_000: DATA = 1'b0;
            15'b10011010_0010_001: DATA = 1'b0;
            15'b10011010_0010_010: DATA = 1'b0;
            15'b10011010_0010_011: DATA = 1'b0;
            15'b10011010_0010_100: DATA = 1'b0;
            15'b10011010_0010_101: DATA = 1'b0;
            15'b10011010_0010_110: DATA = 1'b0;
            15'b10011010_0010_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 1 Row 3
            15'b10011010_0011_000: DATA = 1'b0;
            15'b10011010_0011_001: DATA = 1'b0;
            15'b10011010_0011_010: DATA = 1'b0;
            15'b10011010_0011_011: DATA = 1'b0;
            15'b10011010_0011_100: DATA = 1'b0;
            15'b10011010_0011_101: DATA = 1'b0;
            15'b10011010_0011_110: DATA = 1'b0;
            15'b10011010_0011_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 1 Row 4
            15'b10011010_0100_000: DATA = 1'b0;
            15'b10011010_0100_001: DATA = 1'b0;
            15'b10011010_0100_010: DATA = 1'b0;
            15'b10011010_0100_011: DATA = 1'b0;
            15'b10011010_0100_100: DATA = 1'b0;
            15'b10011010_0100_101: DATA = 1'b0;
            15'b10011010_0100_110: DATA = 1'b0;
            15'b10011010_0100_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 1 Row 5
            15'b10011010_0101_000: DATA = 1'b0;
            15'b10011010_0101_001: DATA = 1'b0;
            15'b10011010_0101_010: DATA = 1'b0;
            15'b10011010_0101_011: DATA = 1'b0;
            15'b10011010_0101_100: DATA = 1'b0;
            15'b10011010_0101_101: DATA = 1'b0;
            15'b10011010_0101_110: DATA = 1'b0;
            15'b10011010_0101_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 1 Row 6
            15'b10011010_0110_000: DATA = 1'b0;
            15'b10011010_0110_001: DATA = 1'b0;
            15'b10011010_0110_010: DATA = 1'b0;
            15'b10011010_0110_011: DATA = 1'b0;
            15'b10011010_0110_100: DATA = 1'b0;
            15'b10011010_0110_101: DATA = 1'b0;
            15'b10011010_0110_110: DATA = 1'b0;
            15'b10011010_0110_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 1 Row 7
            15'b10011010_0111_000: DATA = 1'b0;
            15'b10011010_0111_001: DATA = 1'b0;
            15'b10011010_0111_010: DATA = 1'b0;
            15'b10011010_0111_011: DATA = 1'b0;
            15'b10011010_0111_100: DATA = 1'b0;
            15'b10011010_0111_101: DATA = 1'b0;
            15'b10011010_0111_110: DATA = 1'b0;
            15'b10011010_0111_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 1 Row 8
            15'b10011010_1000_000: DATA = 1'b0;
            15'b10011010_1000_001: DATA = 1'b0;
            15'b10011010_1000_010: DATA = 1'b0;
            15'b10011010_1000_011: DATA = 1'b0;
            15'b10011010_1000_100: DATA = 1'b0;
            15'b10011010_1000_101: DATA = 1'b0;
            15'b10011010_1000_110: DATA = 1'b0;
            15'b10011010_1000_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 1 Row 9
            15'b10011010_1001_000: DATA = 1'b0;
            15'b10011010_1001_001: DATA = 1'b0;
            15'b10011010_1001_010: DATA = 1'b0;
            15'b10011010_1001_011: DATA = 1'b0;
            15'b10011010_1001_100: DATA = 1'b0;
            15'b10011010_1001_101: DATA = 1'b0;
            15'b10011010_1001_110: DATA = 1'b0;
            15'b10011010_1001_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 1 Row 10
            15'b10011010_1010_000: DATA = 1'b0;
            15'b10011010_1010_001: DATA = 1'b0;
            15'b10011010_1010_010: DATA = 1'b0;
            15'b10011010_1010_011: DATA = 1'b0;
            15'b10011010_1010_100: DATA = 1'b0;
            15'b10011010_1010_101: DATA = 1'b0;
            15'b10011010_1010_110: DATA = 1'b0;
            15'b10011010_1010_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 1 Row 11
            15'b10011010_1011_000: DATA = 1'b0;
            15'b10011010_1011_001: DATA = 1'b0;
            15'b10011010_1011_010: DATA = 1'b0;
            15'b10011010_1011_011: DATA = 1'b0;
            15'b10011010_1011_100: DATA = 1'b0;
            15'b10011010_1011_101: DATA = 1'b0;
            15'b10011010_1011_110: DATA = 1'b0;
            15'b10011010_1011_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 1 Row 12
            15'b10011010_1100_000: DATA = 1'b0;
            15'b10011010_1100_001: DATA = 1'b0;
            15'b10011010_1100_010: DATA = 1'b0;
            15'b10011010_1100_011: DATA = 1'b0;
            15'b10011010_1100_100: DATA = 1'b0;
            15'b10011010_1100_101: DATA = 1'b0;
            15'b10011010_1100_110: DATA = 1'b0;
            15'b10011010_1100_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 1 Row 13
            15'b10011010_1101_000: DATA = 1'b0;
            15'b10011010_1101_001: DATA = 1'b0;
            15'b10011010_1101_010: DATA = 1'b0;
            15'b10011010_1101_011: DATA = 1'b0;
            15'b10011010_1101_100: DATA = 1'b0;
            15'b10011010_1101_101: DATA = 1'b0;
            15'b10011010_1101_110: DATA = 1'b0;
            15'b10011010_1101_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 1 Row 14
            15'b10011010_1110_000: DATA = 1'b0;
            15'b10011010_1110_001: DATA = 1'b0;
            15'b10011010_1110_010: DATA = 1'b0;
            15'b10011010_1110_011: DATA = 1'b0;
            15'b10011010_1110_100: DATA = 1'b0;
            15'b10011010_1110_101: DATA = 1'b0;
            15'b10011010_1110_110: DATA = 1'b0;
            15'b10011010_1110_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 1 Row 15
            15'b10011010_1111_000: DATA = 1'b0;
            15'b10011010_1111_001: DATA = 1'b0;
            15'b10011010_1111_010: DATA = 1'b0;
            15'b10011010_1111_011: DATA = 1'b0;
            15'b10011010_1111_100: DATA = 1'b0;
            15'b10011010_1111_101: DATA = 1'b0;
            15'b10011010_1111_110: DATA = 1'b0;
            15'b10011010_1111_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 2 Row 0
            15'b10011011_0000_000: DATA = 1'b0;
            15'b10011011_0000_001: DATA = 1'b0;
            15'b10011011_0000_010: DATA = 1'b0;
            15'b10011011_0000_011: DATA = 1'b0;
            15'b10011011_0000_100: DATA = 1'b0;
            15'b10011011_0000_101: DATA = 1'b0;
            15'b10011011_0000_110: DATA = 1'b0;
            15'b10011011_0000_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 2 Row 1
            15'b10011011_0001_000: DATA = 1'b0;
            15'b10011011_0001_001: DATA = 1'b0;
            15'b10011011_0001_010: DATA = 1'b0;
            15'b10011011_0001_011: DATA = 1'b0;
            15'b10011011_0001_100: DATA = 1'b0;
            15'b10011011_0001_101: DATA = 1'b0;
            15'b10011011_0001_110: DATA = 1'b0;
            15'b10011011_0001_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 2 Row 2
            15'b10011011_0010_000: DATA = 1'b0;
            15'b10011011_0010_001: DATA = 1'b0;
            15'b10011011_0010_010: DATA = 1'b0;
            15'b10011011_0010_011: DATA = 1'b0;
            15'b10011011_0010_100: DATA = 1'b0;
            15'b10011011_0010_101: DATA = 1'b0;
            15'b10011011_0010_110: DATA = 1'b0;
            15'b10011011_0010_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 2 Row 3
            15'b10011011_0011_000: DATA = 1'b0;
            15'b10011011_0011_001: DATA = 1'b0;
            15'b10011011_0011_010: DATA = 1'b0;
            15'b10011011_0011_011: DATA = 1'b0;
            15'b10011011_0011_100: DATA = 1'b0;
            15'b10011011_0011_101: DATA = 1'b0;
            15'b10011011_0011_110: DATA = 1'b0;
            15'b10011011_0011_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 2 Row 4
            15'b10011011_0100_000: DATA = 1'b0;
            15'b10011011_0100_001: DATA = 1'b0;
            15'b10011011_0100_010: DATA = 1'b0;
            15'b10011011_0100_011: DATA = 1'b0;
            15'b10011011_0100_100: DATA = 1'b0;
            15'b10011011_0100_101: DATA = 1'b0;
            15'b10011011_0100_110: DATA = 1'b0;
            15'b10011011_0100_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 2 Row 5
            15'b10011011_0101_000: DATA = 1'b0;
            15'b10011011_0101_001: DATA = 1'b0;
            15'b10011011_0101_010: DATA = 1'b0;
            15'b10011011_0101_011: DATA = 1'b0;
            15'b10011011_0101_100: DATA = 1'b0;
            15'b10011011_0101_101: DATA = 1'b0;
            15'b10011011_0101_110: DATA = 1'b0;
            15'b10011011_0101_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 2 Row 6
            15'b10011011_0110_000: DATA = 1'b0;
            15'b10011011_0110_001: DATA = 1'b0;
            15'b10011011_0110_010: DATA = 1'b0;
            15'b10011011_0110_011: DATA = 1'b0;
            15'b10011011_0110_100: DATA = 1'b0;
            15'b10011011_0110_101: DATA = 1'b0;
            15'b10011011_0110_110: DATA = 1'b0;
            15'b10011011_0110_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 2 Row 7
            15'b10011011_0111_000: DATA = 1'b0;
            15'b10011011_0111_001: DATA = 1'b0;
            15'b10011011_0111_010: DATA = 1'b0;
            15'b10011011_0111_011: DATA = 1'b0;
            15'b10011011_0111_100: DATA = 1'b0;
            15'b10011011_0111_101: DATA = 1'b0;
            15'b10011011_0111_110: DATA = 1'b0;
            15'b10011011_0111_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 2 Row 8
            15'b10011011_1000_000: DATA = 1'b0;
            15'b10011011_1000_001: DATA = 1'b0;
            15'b10011011_1000_010: DATA = 1'b0;
            15'b10011011_1000_011: DATA = 1'b0;
            15'b10011011_1000_100: DATA = 1'b0;
            15'b10011011_1000_101: DATA = 1'b0;
            15'b10011011_1000_110: DATA = 1'b0;
            15'b10011011_1000_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 2 Row 9
            15'b10011011_1001_000: DATA = 1'b0;
            15'b10011011_1001_001: DATA = 1'b0;
            15'b10011011_1001_010: DATA = 1'b0;
            15'b10011011_1001_011: DATA = 1'b0;
            15'b10011011_1001_100: DATA = 1'b0;
            15'b10011011_1001_101: DATA = 1'b0;
            15'b10011011_1001_110: DATA = 1'b0;
            15'b10011011_1001_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 2 Row 10
            15'b10011011_1010_000: DATA = 1'b0;
            15'b10011011_1010_001: DATA = 1'b0;
            15'b10011011_1010_010: DATA = 1'b0;
            15'b10011011_1010_011: DATA = 1'b0;
            15'b10011011_1010_100: DATA = 1'b0;
            15'b10011011_1010_101: DATA = 1'b0;
            15'b10011011_1010_110: DATA = 1'b0;
            15'b10011011_1010_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 2 Row 11
            15'b10011011_1011_000: DATA = 1'b0;
            15'b10011011_1011_001: DATA = 1'b0;
            15'b10011011_1011_010: DATA = 1'b0;
            15'b10011011_1011_011: DATA = 1'b0;
            15'b10011011_1011_100: DATA = 1'b0;
            15'b10011011_1011_101: DATA = 1'b0;
            15'b10011011_1011_110: DATA = 1'b0;
            15'b10011011_1011_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 2 Row 12
            15'b10011011_1100_000: DATA = 1'b0;
            15'b10011011_1100_001: DATA = 1'b0;
            15'b10011011_1100_010: DATA = 1'b0;
            15'b10011011_1100_011: DATA = 1'b0;
            15'b10011011_1100_100: DATA = 1'b0;
            15'b10011011_1100_101: DATA = 1'b0;
            15'b10011011_1100_110: DATA = 1'b0;
            15'b10011011_1100_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 2 Row 13
            15'b10011011_1101_000: DATA = 1'b0;
            15'b10011011_1101_001: DATA = 1'b0;
            15'b10011011_1101_010: DATA = 1'b0;
            15'b10011011_1101_011: DATA = 1'b0;
            15'b10011011_1101_100: DATA = 1'b0;
            15'b10011011_1101_101: DATA = 1'b0;
            15'b10011011_1101_110: DATA = 1'b0;
            15'b10011011_1101_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 2 Row 14
            15'b10011011_1110_000: DATA = 1'b0;
            15'b10011011_1110_001: DATA = 1'b0;
            15'b10011011_1110_010: DATA = 1'b0;
            15'b10011011_1110_011: DATA = 1'b0;
            15'b10011011_1110_100: DATA = 1'b0;
            15'b10011011_1110_101: DATA = 1'b0;
            15'b10011011_1110_110: DATA = 1'b0;
            15'b10011011_1110_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 2 Row 15
            15'b10011011_1111_000: DATA = 1'b0;
            15'b10011011_1111_001: DATA = 1'b0;
            15'b10011011_1111_010: DATA = 1'b0;
            15'b10011011_1111_011: DATA = 1'b0;
            15'b10011011_1111_100: DATA = 1'b0;
            15'b10011011_1111_101: DATA = 1'b0;
            15'b10011011_1111_110: DATA = 1'b0;
            15'b10011011_1111_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 3 Row 0
            15'b10011100_0000_000: DATA = 1'b0;
            15'b10011100_0000_001: DATA = 1'b0;
            15'b10011100_0000_010: DATA = 1'b0;
            15'b10011100_0000_011: DATA = 1'b0;
            15'b10011100_0000_100: DATA = 1'b0;
            15'b10011100_0000_101: DATA = 1'b0;
            15'b10011100_0000_110: DATA = 1'b0;
            15'b10011100_0000_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 3 Row 1
            15'b10011100_0001_000: DATA = 1'b0;
            15'b10011100_0001_001: DATA = 1'b0;
            15'b10011100_0001_010: DATA = 1'b0;
            15'b10011100_0001_011: DATA = 1'b0;
            15'b10011100_0001_100: DATA = 1'b0;
            15'b10011100_0001_101: DATA = 1'b0;
            15'b10011100_0001_110: DATA = 1'b0;
            15'b10011100_0001_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 3 Row 2
            15'b10011100_0010_000: DATA = 1'b0;
            15'b10011100_0010_001: DATA = 1'b0;
            15'b10011100_0010_010: DATA = 1'b0;
            15'b10011100_0010_011: DATA = 1'b0;
            15'b10011100_0010_100: DATA = 1'b0;
            15'b10011100_0010_101: DATA = 1'b0;
            15'b10011100_0010_110: DATA = 1'b0;
            15'b10011100_0010_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 3 Row 3
            15'b10011100_0011_000: DATA = 1'b0;
            15'b10011100_0011_001: DATA = 1'b0;
            15'b10011100_0011_010: DATA = 1'b0;
            15'b10011100_0011_011: DATA = 1'b0;
            15'b10011100_0011_100: DATA = 1'b0;
            15'b10011100_0011_101: DATA = 1'b0;
            15'b10011100_0011_110: DATA = 1'b0;
            15'b10011100_0011_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 3 Row 4
            15'b10011100_0100_000: DATA = 1'b0;
            15'b10011100_0100_001: DATA = 1'b0;
            15'b10011100_0100_010: DATA = 1'b0;
            15'b10011100_0100_011: DATA = 1'b0;
            15'b10011100_0100_100: DATA = 1'b0;
            15'b10011100_0100_101: DATA = 1'b0;
            15'b10011100_0100_110: DATA = 1'b0;
            15'b10011100_0100_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 3 Row 5
            15'b10011100_0101_000: DATA = 1'b0;
            15'b10011100_0101_001: DATA = 1'b0;
            15'b10011100_0101_010: DATA = 1'b0;
            15'b10011100_0101_011: DATA = 1'b0;
            15'b10011100_0101_100: DATA = 1'b0;
            15'b10011100_0101_101: DATA = 1'b0;
            15'b10011100_0101_110: DATA = 1'b0;
            15'b10011100_0101_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 3 Row 6
            15'b10011100_0110_000: DATA = 1'b0;
            15'b10011100_0110_001: DATA = 1'b0;
            15'b10011100_0110_010: DATA = 1'b0;
            15'b10011100_0110_011: DATA = 1'b0;
            15'b10011100_0110_100: DATA = 1'b0;
            15'b10011100_0110_101: DATA = 1'b0;
            15'b10011100_0110_110: DATA = 1'b0;
            15'b10011100_0110_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 3 Row 7
            15'b10011100_0111_000: DATA = 1'b0;
            15'b10011100_0111_001: DATA = 1'b0;
            15'b10011100_0111_010: DATA = 1'b0;
            15'b10011100_0111_011: DATA = 1'b0;
            15'b10011100_0111_100: DATA = 1'b0;
            15'b10011100_0111_101: DATA = 1'b0;
            15'b10011100_0111_110: DATA = 1'b0;
            15'b10011100_0111_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 3 Row 8
            15'b10011100_1000_000: DATA = 1'b0;
            15'b10011100_1000_001: DATA = 1'b0;
            15'b10011100_1000_010: DATA = 1'b0;
            15'b10011100_1000_011: DATA = 1'b0;
            15'b10011100_1000_100: DATA = 1'b0;
            15'b10011100_1000_101: DATA = 1'b0;
            15'b10011100_1000_110: DATA = 1'b0;
            15'b10011100_1000_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 3 Row 9
            15'b10011100_1001_000: DATA = 1'b0;
            15'b10011100_1001_001: DATA = 1'b0;
            15'b10011100_1001_010: DATA = 1'b0;
            15'b10011100_1001_011: DATA = 1'b0;
            15'b10011100_1001_100: DATA = 1'b0;
            15'b10011100_1001_101: DATA = 1'b0;
            15'b10011100_1001_110: DATA = 1'b0;
            15'b10011100_1001_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 3 Row 10
            15'b10011100_1010_000: DATA = 1'b0;
            15'b10011100_1010_001: DATA = 1'b0;
            15'b10011100_1010_010: DATA = 1'b0;
            15'b10011100_1010_011: DATA = 1'b0;
            15'b10011100_1010_100: DATA = 1'b0;
            15'b10011100_1010_101: DATA = 1'b0;
            15'b10011100_1010_110: DATA = 1'b0;
            15'b10011100_1010_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 3 Row 11
            15'b10011100_1011_000: DATA = 1'b0;
            15'b10011100_1011_001: DATA = 1'b0;
            15'b10011100_1011_010: DATA = 1'b0;
            15'b10011100_1011_011: DATA = 1'b0;
            15'b10011100_1011_100: DATA = 1'b0;
            15'b10011100_1011_101: DATA = 1'b0;
            15'b10011100_1011_110: DATA = 1'b0;
            15'b10011100_1011_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 3 Row 12
            15'b10011100_1100_000: DATA = 1'b0;
            15'b10011100_1100_001: DATA = 1'b0;
            15'b10011100_1100_010: DATA = 1'b0;
            15'b10011100_1100_011: DATA = 1'b0;
            15'b10011100_1100_100: DATA = 1'b0;
            15'b10011100_1100_101: DATA = 1'b0;
            15'b10011100_1100_110: DATA = 1'b0;
            15'b10011100_1100_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 3 Row 13
            15'b10011100_1101_000: DATA = 1'b0;
            15'b10011100_1101_001: DATA = 1'b0;
            15'b10011100_1101_010: DATA = 1'b0;
            15'b10011100_1101_011: DATA = 1'b0;
            15'b10011100_1101_100: DATA = 1'b0;
            15'b10011100_1101_101: DATA = 1'b0;
            15'b10011100_1101_110: DATA = 1'b0;
            15'b10011100_1101_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 3 Row 14
            15'b10011100_1110_000: DATA = 1'b0;
            15'b10011100_1110_001: DATA = 1'b0;
            15'b10011100_1110_010: DATA = 1'b0;
            15'b10011100_1110_011: DATA = 1'b0;
            15'b10011100_1110_100: DATA = 1'b0;
            15'b10011100_1110_101: DATA = 1'b0;
            15'b10011100_1110_110: DATA = 1'b0;
            15'b10011100_1110_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 3 Row 15
            15'b10011100_1111_000: DATA = 1'b0;
            15'b10011100_1111_001: DATA = 1'b0;
            15'b10011100_1111_010: DATA = 1'b0;
            15'b10011100_1111_011: DATA = 1'b0;
            15'b10011100_1111_100: DATA = 1'b0;
            15'b10011100_1111_101: DATA = 1'b0;
            15'b10011100_1111_110: DATA = 1'b0;
            15'b10011100_1111_111: DATA = 1'b0;
            // SQUARE+ ROW 1 COL 4 Row 0
            15'b10011101_0000_000: DATA = 1'b0;
            15'b10011101_0000_001: DATA = 1'b0;
            15'b10011101_0000_010: DATA = 1'b0;
            15'b10011101_0000_011: DATA = 1'b0;
            15'b10011101_0000_100: DATA = 1'b0;
            15'b10011101_0000_101: DATA = 1'b0;
            15'b10011101_0000_110: DATA = 1'b0;
            15'b10011101_0000_111: DATA = 1'b1;
            // SQUARE+ ROW 1 COL 4 Row 1
            15'b10011101_0001_000: DATA = 1'b0;
            15'b10011101_0001_001: DATA = 1'b0;
            15'b10011101_0001_010: DATA = 1'b0;
            15'b10011101_0001_011: DATA = 1'b0;
            15'b10011101_0001_100: DATA = 1'b0;
            15'b10011101_0001_101: DATA = 1'b0;
            15'b10011101_0001_110: DATA = 1'b0;
            15'b10011101_0001_111: DATA = 1'b1;
            // SQUARE+ ROW 1 COL 4 Row 2
            15'b10011101_0010_000: DATA = 1'b0;
            15'b10011101_0010_001: DATA = 1'b0;
            15'b10011101_0010_010: DATA = 1'b0;
            15'b10011101_0010_011: DATA = 1'b0;
            15'b10011101_0010_100: DATA = 1'b0;
            15'b10011101_0010_101: DATA = 1'b0;
            15'b10011101_0010_110: DATA = 1'b0;
            15'b10011101_0010_111: DATA = 1'b1;
            // SQUARE+ ROW 1 COL 4 Row 3
            15'b10011101_0011_000: DATA = 1'b0;
            15'b10011101_0011_001: DATA = 1'b0;
            15'b10011101_0011_010: DATA = 1'b0;
            15'b10011101_0011_011: DATA = 1'b0;
            15'b10011101_0011_100: DATA = 1'b0;
            15'b10011101_0011_101: DATA = 1'b0;
            15'b10011101_0011_110: DATA = 1'b0;
            15'b10011101_0011_111: DATA = 1'b1;
            // SQUARE+ ROW 1 COL 4 Row 4
            15'b10011101_0100_000: DATA = 1'b0;
            15'b10011101_0100_001: DATA = 1'b0;
            15'b10011101_0100_010: DATA = 1'b0;
            15'b10011101_0100_011: DATA = 1'b0;
            15'b10011101_0100_100: DATA = 1'b0;
            15'b10011101_0100_101: DATA = 1'b0;
            15'b10011101_0100_110: DATA = 1'b0;
            15'b10011101_0100_111: DATA = 1'b1;
            // SQUARE+ ROW 1 COL 4 Row 5
            15'b10011101_0101_000: DATA = 1'b0;
            15'b10011101_0101_001: DATA = 1'b0;
            15'b10011101_0101_010: DATA = 1'b0;
            15'b10011101_0101_011: DATA = 1'b0;
            15'b10011101_0101_100: DATA = 1'b0;
            15'b10011101_0101_101: DATA = 1'b0;
            15'b10011101_0101_110: DATA = 1'b0;
            15'b10011101_0101_111: DATA = 1'b1;
            // SQUARE+ ROW 1 COL 4 Row 6
            15'b10011101_0110_000: DATA = 1'b0;
            15'b10011101_0110_001: DATA = 1'b0;
            15'b10011101_0110_010: DATA = 1'b0;
            15'b10011101_0110_011: DATA = 1'b0;
            15'b10011101_0110_100: DATA = 1'b0;
            15'b10011101_0110_101: DATA = 1'b0;
            15'b10011101_0110_110: DATA = 1'b0;
            15'b10011101_0110_111: DATA = 1'b1;
            // SQUARE+ ROW 1 COL 4 Row 7
            15'b10011101_0111_000: DATA = 1'b0;
            15'b10011101_0111_001: DATA = 1'b0;
            15'b10011101_0111_010: DATA = 1'b0;
            15'b10011101_0111_011: DATA = 1'b0;
            15'b10011101_0111_100: DATA = 1'b0;
            15'b10011101_0111_101: DATA = 1'b0;
            15'b10011101_0111_110: DATA = 1'b0;
            15'b10011101_0111_111: DATA = 1'b1;
            // SQUARE+ ROW 1 COL 4 Row 8
            15'b10011101_1000_000: DATA = 1'b0;
            15'b10011101_1000_001: DATA = 1'b0;
            15'b10011101_1000_010: DATA = 1'b0;
            15'b10011101_1000_011: DATA = 1'b0;
            15'b10011101_1000_100: DATA = 1'b0;
            15'b10011101_1000_101: DATA = 1'b0;
            15'b10011101_1000_110: DATA = 1'b0;
            15'b10011101_1000_111: DATA = 1'b1;
            // SQUARE+ ROW 1 COL 4 Row 9
            15'b10011101_1001_000: DATA = 1'b0;
            15'b10011101_1001_001: DATA = 1'b0;
            15'b10011101_1001_010: DATA = 1'b0;
            15'b10011101_1001_011: DATA = 1'b0;
            15'b10011101_1001_100: DATA = 1'b0;
            15'b10011101_1001_101: DATA = 1'b0;
            15'b10011101_1001_110: DATA = 1'b0;
            15'b10011101_1001_111: DATA = 1'b1;
            // SQUARE+ ROW 1 COL 4 Row 10
            15'b10011101_1010_000: DATA = 1'b0;
            15'b10011101_1010_001: DATA = 1'b0;
            15'b10011101_1010_010: DATA = 1'b0;
            15'b10011101_1010_011: DATA = 1'b0;
            15'b10011101_1010_100: DATA = 1'b0;
            15'b10011101_1010_101: DATA = 1'b0;
            15'b10011101_1010_110: DATA = 1'b0;
            15'b10011101_1010_111: DATA = 1'b1;
            // SQUARE+ ROW 1 COL 4 Row 11
            15'b10011101_1011_000: DATA = 1'b0;
            15'b10011101_1011_001: DATA = 1'b0;
            15'b10011101_1011_010: DATA = 1'b0;
            15'b10011101_1011_011: DATA = 1'b0;
            15'b10011101_1011_100: DATA = 1'b0;
            15'b10011101_1011_101: DATA = 1'b0;
            15'b10011101_1011_110: DATA = 1'b0;
            15'b10011101_1011_111: DATA = 1'b1;
            // SQUARE+ ROW 1 COL 4 Row 12
            15'b10011101_1100_000: DATA = 1'b0;
            15'b10011101_1100_001: DATA = 1'b0;
            15'b10011101_1100_010: DATA = 1'b0;
            15'b10011101_1100_011: DATA = 1'b0;
            15'b10011101_1100_100: DATA = 1'b0;
            15'b10011101_1100_101: DATA = 1'b0;
            15'b10011101_1100_110: DATA = 1'b0;
            15'b10011101_1100_111: DATA = 1'b1;
            // SQUARE+ ROW 1 COL 4 Row 13
            15'b10011101_1101_000: DATA = 1'b0;
            15'b10011101_1101_001: DATA = 1'b0;
            15'b10011101_1101_010: DATA = 1'b0;
            15'b10011101_1101_011: DATA = 1'b0;
            15'b10011101_1101_100: DATA = 1'b0;
            15'b10011101_1101_101: DATA = 1'b0;
            15'b10011101_1101_110: DATA = 1'b0;
            15'b10011101_1101_111: DATA = 1'b1;
            // SQUARE+ ROW 1 COL 4 Row 14
            15'b10011101_1110_000: DATA = 1'b0;
            15'b10011101_1110_001: DATA = 1'b0;
            15'b10011101_1110_010: DATA = 1'b0;
            15'b10011101_1110_011: DATA = 1'b0;
            15'b10011101_1110_100: DATA = 1'b0;
            15'b10011101_1110_101: DATA = 1'b0;
            15'b10011101_1110_110: DATA = 1'b0;
            15'b10011101_1110_111: DATA = 1'b1;
            // SQUARE+ ROW 1 COL 4 Row 15
            15'b10011101_1111_000: DATA = 1'b0;
            15'b10011101_1111_001: DATA = 1'b0;
            15'b10011101_1111_010: DATA = 1'b0;
            15'b10011101_1111_011: DATA = 1'b0;
            15'b10011101_1111_100: DATA = 1'b0;
            15'b10011101_1111_101: DATA = 1'b0;
            15'b10011101_1111_110: DATA = 1'b0;
            15'b10011101_1111_111: DATA = 1'b1;
            // SQUARE- ROW 0 COL 0 Row 0
            15'b10011110_0000_000: DATA = 1'b1;
            15'b10011110_0000_001: DATA = 1'b0;
            15'b10011110_0000_010: DATA = 1'b0;
            15'b10011110_0000_011: DATA = 1'b0;
            15'b10011110_0000_100: DATA = 1'b0;
            15'b10011110_0000_101: DATA = 1'b0;
            15'b10011110_0000_110: DATA = 1'b0;
            15'b10011110_0000_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 0 Row 1
            15'b10011110_0001_000: DATA = 1'b1;
            15'b10011110_0001_001: DATA = 1'b0;
            15'b10011110_0001_010: DATA = 1'b0;
            15'b10011110_0001_011: DATA = 1'b0;
            15'b10011110_0001_100: DATA = 1'b0;
            15'b10011110_0001_101: DATA = 1'b0;
            15'b10011110_0001_110: DATA = 1'b0;
            15'b10011110_0001_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 0 Row 2
            15'b10011110_0010_000: DATA = 1'b1;
            15'b10011110_0010_001: DATA = 1'b0;
            15'b10011110_0010_010: DATA = 1'b0;
            15'b10011110_0010_011: DATA = 1'b0;
            15'b10011110_0010_100: DATA = 1'b0;
            15'b10011110_0010_101: DATA = 1'b0;
            15'b10011110_0010_110: DATA = 1'b0;
            15'b10011110_0010_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 0 Row 3
            15'b10011110_0011_000: DATA = 1'b1;
            15'b10011110_0011_001: DATA = 1'b0;
            15'b10011110_0011_010: DATA = 1'b0;
            15'b10011110_0011_011: DATA = 1'b0;
            15'b10011110_0011_100: DATA = 1'b0;
            15'b10011110_0011_101: DATA = 1'b0;
            15'b10011110_0011_110: DATA = 1'b0;
            15'b10011110_0011_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 0 Row 4
            15'b10011110_0100_000: DATA = 1'b1;
            15'b10011110_0100_001: DATA = 1'b0;
            15'b10011110_0100_010: DATA = 1'b0;
            15'b10011110_0100_011: DATA = 1'b0;
            15'b10011110_0100_100: DATA = 1'b0;
            15'b10011110_0100_101: DATA = 1'b0;
            15'b10011110_0100_110: DATA = 1'b0;
            15'b10011110_0100_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 0 Row 5
            15'b10011110_0101_000: DATA = 1'b1;
            15'b10011110_0101_001: DATA = 1'b0;
            15'b10011110_0101_010: DATA = 1'b0;
            15'b10011110_0101_011: DATA = 1'b0;
            15'b10011110_0101_100: DATA = 1'b0;
            15'b10011110_0101_101: DATA = 1'b0;
            15'b10011110_0101_110: DATA = 1'b0;
            15'b10011110_0101_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 0 Row 6
            15'b10011110_0110_000: DATA = 1'b1;
            15'b10011110_0110_001: DATA = 1'b0;
            15'b10011110_0110_010: DATA = 1'b0;
            15'b10011110_0110_011: DATA = 1'b0;
            15'b10011110_0110_100: DATA = 1'b0;
            15'b10011110_0110_101: DATA = 1'b0;
            15'b10011110_0110_110: DATA = 1'b0;
            15'b10011110_0110_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 0 Row 7
            15'b10011110_0111_000: DATA = 1'b1;
            15'b10011110_0111_001: DATA = 1'b0;
            15'b10011110_0111_010: DATA = 1'b0;
            15'b10011110_0111_011: DATA = 1'b0;
            15'b10011110_0111_100: DATA = 1'b0;
            15'b10011110_0111_101: DATA = 1'b0;
            15'b10011110_0111_110: DATA = 1'b0;
            15'b10011110_0111_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 0 Row 8
            15'b10011110_1000_000: DATA = 1'b1;
            15'b10011110_1000_001: DATA = 1'b0;
            15'b10011110_1000_010: DATA = 1'b0;
            15'b10011110_1000_011: DATA = 1'b0;
            15'b10011110_1000_100: DATA = 1'b0;
            15'b10011110_1000_101: DATA = 1'b0;
            15'b10011110_1000_110: DATA = 1'b0;
            15'b10011110_1000_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 0 Row 9
            15'b10011110_1001_000: DATA = 1'b1;
            15'b10011110_1001_001: DATA = 1'b0;
            15'b10011110_1001_010: DATA = 1'b0;
            15'b10011110_1001_011: DATA = 1'b0;
            15'b10011110_1001_100: DATA = 1'b0;
            15'b10011110_1001_101: DATA = 1'b0;
            15'b10011110_1001_110: DATA = 1'b0;
            15'b10011110_1001_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 0 Row 10
            15'b10011110_1010_000: DATA = 1'b1;
            15'b10011110_1010_001: DATA = 1'b0;
            15'b10011110_1010_010: DATA = 1'b0;
            15'b10011110_1010_011: DATA = 1'b0;
            15'b10011110_1010_100: DATA = 1'b0;
            15'b10011110_1010_101: DATA = 1'b0;
            15'b10011110_1010_110: DATA = 1'b0;
            15'b10011110_1010_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 0 Row 11
            15'b10011110_1011_000: DATA = 1'b1;
            15'b10011110_1011_001: DATA = 1'b0;
            15'b10011110_1011_010: DATA = 1'b0;
            15'b10011110_1011_011: DATA = 1'b0;
            15'b10011110_1011_100: DATA = 1'b0;
            15'b10011110_1011_101: DATA = 1'b0;
            15'b10011110_1011_110: DATA = 1'b0;
            15'b10011110_1011_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 0 Row 12
            15'b10011110_1100_000: DATA = 1'b1;
            15'b10011110_1100_001: DATA = 1'b0;
            15'b10011110_1100_010: DATA = 1'b0;
            15'b10011110_1100_011: DATA = 1'b0;
            15'b10011110_1100_100: DATA = 1'b0;
            15'b10011110_1100_101: DATA = 1'b0;
            15'b10011110_1100_110: DATA = 1'b0;
            15'b10011110_1100_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 0 Row 13
            15'b10011110_1101_000: DATA = 1'b1;
            15'b10011110_1101_001: DATA = 1'b0;
            15'b10011110_1101_010: DATA = 1'b0;
            15'b10011110_1101_011: DATA = 1'b0;
            15'b10011110_1101_100: DATA = 1'b0;
            15'b10011110_1101_101: DATA = 1'b0;
            15'b10011110_1101_110: DATA = 1'b0;
            15'b10011110_1101_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 0 Row 14
            15'b10011110_1110_000: DATA = 1'b1;
            15'b10011110_1110_001: DATA = 1'b0;
            15'b10011110_1110_010: DATA = 1'b0;
            15'b10011110_1110_011: DATA = 1'b0;
            15'b10011110_1110_100: DATA = 1'b0;
            15'b10011110_1110_101: DATA = 1'b0;
            15'b10011110_1110_110: DATA = 1'b0;
            15'b10011110_1110_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 0 Row 15
            15'b10011110_1111_000: DATA = 1'b1;
            15'b10011110_1111_001: DATA = 1'b0;
            15'b10011110_1111_010: DATA = 1'b0;
            15'b10011110_1111_011: DATA = 1'b0;
            15'b10011110_1111_100: DATA = 1'b0;
            15'b10011110_1111_101: DATA = 1'b0;
            15'b10011110_1111_110: DATA = 1'b0;
            15'b10011110_1111_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 1 Row 0
            15'b10011111_0000_000: DATA = 1'b0;
            15'b10011111_0000_001: DATA = 1'b0;
            15'b10011111_0000_010: DATA = 1'b0;
            15'b10011111_0000_011: DATA = 1'b0;
            15'b10011111_0000_100: DATA = 1'b0;
            15'b10011111_0000_101: DATA = 1'b0;
            15'b10011111_0000_110: DATA = 1'b0;
            15'b10011111_0000_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 1 Row 1
            15'b10011111_0001_000: DATA = 1'b0;
            15'b10011111_0001_001: DATA = 1'b0;
            15'b10011111_0001_010: DATA = 1'b0;
            15'b10011111_0001_011: DATA = 1'b0;
            15'b10011111_0001_100: DATA = 1'b0;
            15'b10011111_0001_101: DATA = 1'b0;
            15'b10011111_0001_110: DATA = 1'b0;
            15'b10011111_0001_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 1 Row 2
            15'b10011111_0010_000: DATA = 1'b0;
            15'b10011111_0010_001: DATA = 1'b0;
            15'b10011111_0010_010: DATA = 1'b0;
            15'b10011111_0010_011: DATA = 1'b0;
            15'b10011111_0010_100: DATA = 1'b0;
            15'b10011111_0010_101: DATA = 1'b0;
            15'b10011111_0010_110: DATA = 1'b0;
            15'b10011111_0010_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 1 Row 3
            15'b10011111_0011_000: DATA = 1'b0;
            15'b10011111_0011_001: DATA = 1'b0;
            15'b10011111_0011_010: DATA = 1'b0;
            15'b10011111_0011_011: DATA = 1'b0;
            15'b10011111_0011_100: DATA = 1'b0;
            15'b10011111_0011_101: DATA = 1'b0;
            15'b10011111_0011_110: DATA = 1'b0;
            15'b10011111_0011_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 1 Row 4
            15'b10011111_0100_000: DATA = 1'b0;
            15'b10011111_0100_001: DATA = 1'b0;
            15'b10011111_0100_010: DATA = 1'b0;
            15'b10011111_0100_011: DATA = 1'b0;
            15'b10011111_0100_100: DATA = 1'b0;
            15'b10011111_0100_101: DATA = 1'b0;
            15'b10011111_0100_110: DATA = 1'b0;
            15'b10011111_0100_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 1 Row 5
            15'b10011111_0101_000: DATA = 1'b0;
            15'b10011111_0101_001: DATA = 1'b0;
            15'b10011111_0101_010: DATA = 1'b0;
            15'b10011111_0101_011: DATA = 1'b0;
            15'b10011111_0101_100: DATA = 1'b0;
            15'b10011111_0101_101: DATA = 1'b0;
            15'b10011111_0101_110: DATA = 1'b0;
            15'b10011111_0101_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 1 Row 6
            15'b10011111_0110_000: DATA = 1'b0;
            15'b10011111_0110_001: DATA = 1'b0;
            15'b10011111_0110_010: DATA = 1'b0;
            15'b10011111_0110_011: DATA = 1'b0;
            15'b10011111_0110_100: DATA = 1'b0;
            15'b10011111_0110_101: DATA = 1'b0;
            15'b10011111_0110_110: DATA = 1'b0;
            15'b10011111_0110_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 1 Row 7
            15'b10011111_0111_000: DATA = 1'b0;
            15'b10011111_0111_001: DATA = 1'b0;
            15'b10011111_0111_010: DATA = 1'b0;
            15'b10011111_0111_011: DATA = 1'b0;
            15'b10011111_0111_100: DATA = 1'b0;
            15'b10011111_0111_101: DATA = 1'b0;
            15'b10011111_0111_110: DATA = 1'b0;
            15'b10011111_0111_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 1 Row 8
            15'b10011111_1000_000: DATA = 1'b0;
            15'b10011111_1000_001: DATA = 1'b0;
            15'b10011111_1000_010: DATA = 1'b0;
            15'b10011111_1000_011: DATA = 1'b0;
            15'b10011111_1000_100: DATA = 1'b0;
            15'b10011111_1000_101: DATA = 1'b0;
            15'b10011111_1000_110: DATA = 1'b0;
            15'b10011111_1000_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 1 Row 9
            15'b10011111_1001_000: DATA = 1'b0;
            15'b10011111_1001_001: DATA = 1'b0;
            15'b10011111_1001_010: DATA = 1'b0;
            15'b10011111_1001_011: DATA = 1'b0;
            15'b10011111_1001_100: DATA = 1'b0;
            15'b10011111_1001_101: DATA = 1'b0;
            15'b10011111_1001_110: DATA = 1'b0;
            15'b10011111_1001_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 1 Row 10
            15'b10011111_1010_000: DATA = 1'b0;
            15'b10011111_1010_001: DATA = 1'b0;
            15'b10011111_1010_010: DATA = 1'b0;
            15'b10011111_1010_011: DATA = 1'b0;
            15'b10011111_1010_100: DATA = 1'b0;
            15'b10011111_1010_101: DATA = 1'b0;
            15'b10011111_1010_110: DATA = 1'b0;
            15'b10011111_1010_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 1 Row 11
            15'b10011111_1011_000: DATA = 1'b0;
            15'b10011111_1011_001: DATA = 1'b0;
            15'b10011111_1011_010: DATA = 1'b0;
            15'b10011111_1011_011: DATA = 1'b0;
            15'b10011111_1011_100: DATA = 1'b0;
            15'b10011111_1011_101: DATA = 1'b0;
            15'b10011111_1011_110: DATA = 1'b0;
            15'b10011111_1011_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 1 Row 12
            15'b10011111_1100_000: DATA = 1'b0;
            15'b10011111_1100_001: DATA = 1'b0;
            15'b10011111_1100_010: DATA = 1'b0;
            15'b10011111_1100_011: DATA = 1'b0;
            15'b10011111_1100_100: DATA = 1'b0;
            15'b10011111_1100_101: DATA = 1'b0;
            15'b10011111_1100_110: DATA = 1'b0;
            15'b10011111_1100_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 1 Row 13
            15'b10011111_1101_000: DATA = 1'b0;
            15'b10011111_1101_001: DATA = 1'b0;
            15'b10011111_1101_010: DATA = 1'b0;
            15'b10011111_1101_011: DATA = 1'b0;
            15'b10011111_1101_100: DATA = 1'b0;
            15'b10011111_1101_101: DATA = 1'b0;
            15'b10011111_1101_110: DATA = 1'b0;
            15'b10011111_1101_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 1 Row 14
            15'b10011111_1110_000: DATA = 1'b0;
            15'b10011111_1110_001: DATA = 1'b0;
            15'b10011111_1110_010: DATA = 1'b0;
            15'b10011111_1110_011: DATA = 1'b0;
            15'b10011111_1110_100: DATA = 1'b0;
            15'b10011111_1110_101: DATA = 1'b0;
            15'b10011111_1110_110: DATA = 1'b0;
            15'b10011111_1110_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 1 Row 15
            15'b10011111_1111_000: DATA = 1'b0;
            15'b10011111_1111_001: DATA = 1'b0;
            15'b10011111_1111_010: DATA = 1'b0;
            15'b10011111_1111_011: DATA = 1'b0;
            15'b10011111_1111_100: DATA = 1'b0;
            15'b10011111_1111_101: DATA = 1'b0;
            15'b10011111_1111_110: DATA = 1'b0;
            15'b10011111_1111_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 2 Row 0
            15'b10100000_0000_000: DATA = 1'b0;
            15'b10100000_0000_001: DATA = 1'b0;
            15'b10100000_0000_010: DATA = 1'b0;
            15'b10100000_0000_011: DATA = 1'b0;
            15'b10100000_0000_100: DATA = 1'b0;
            15'b10100000_0000_101: DATA = 1'b0;
            15'b10100000_0000_110: DATA = 1'b0;
            15'b10100000_0000_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 2 Row 1
            15'b10100000_0001_000: DATA = 1'b0;
            15'b10100000_0001_001: DATA = 1'b0;
            15'b10100000_0001_010: DATA = 1'b0;
            15'b10100000_0001_011: DATA = 1'b0;
            15'b10100000_0001_100: DATA = 1'b0;
            15'b10100000_0001_101: DATA = 1'b0;
            15'b10100000_0001_110: DATA = 1'b0;
            15'b10100000_0001_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 2 Row 2
            15'b10100000_0010_000: DATA = 1'b0;
            15'b10100000_0010_001: DATA = 1'b0;
            15'b10100000_0010_010: DATA = 1'b0;
            15'b10100000_0010_011: DATA = 1'b0;
            15'b10100000_0010_100: DATA = 1'b0;
            15'b10100000_0010_101: DATA = 1'b0;
            15'b10100000_0010_110: DATA = 1'b0;
            15'b10100000_0010_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 2 Row 3
            15'b10100000_0011_000: DATA = 1'b0;
            15'b10100000_0011_001: DATA = 1'b0;
            15'b10100000_0011_010: DATA = 1'b0;
            15'b10100000_0011_011: DATA = 1'b0;
            15'b10100000_0011_100: DATA = 1'b0;
            15'b10100000_0011_101: DATA = 1'b0;
            15'b10100000_0011_110: DATA = 1'b0;
            15'b10100000_0011_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 2 Row 4
            15'b10100000_0100_000: DATA = 1'b0;
            15'b10100000_0100_001: DATA = 1'b0;
            15'b10100000_0100_010: DATA = 1'b0;
            15'b10100000_0100_011: DATA = 1'b0;
            15'b10100000_0100_100: DATA = 1'b0;
            15'b10100000_0100_101: DATA = 1'b0;
            15'b10100000_0100_110: DATA = 1'b0;
            15'b10100000_0100_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 2 Row 5
            15'b10100000_0101_000: DATA = 1'b0;
            15'b10100000_0101_001: DATA = 1'b0;
            15'b10100000_0101_010: DATA = 1'b0;
            15'b10100000_0101_011: DATA = 1'b0;
            15'b10100000_0101_100: DATA = 1'b0;
            15'b10100000_0101_101: DATA = 1'b0;
            15'b10100000_0101_110: DATA = 1'b0;
            15'b10100000_0101_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 2 Row 6
            15'b10100000_0110_000: DATA = 1'b0;
            15'b10100000_0110_001: DATA = 1'b0;
            15'b10100000_0110_010: DATA = 1'b0;
            15'b10100000_0110_011: DATA = 1'b0;
            15'b10100000_0110_100: DATA = 1'b0;
            15'b10100000_0110_101: DATA = 1'b0;
            15'b10100000_0110_110: DATA = 1'b0;
            15'b10100000_0110_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 2 Row 7
            15'b10100000_0111_000: DATA = 1'b0;
            15'b10100000_0111_001: DATA = 1'b0;
            15'b10100000_0111_010: DATA = 1'b0;
            15'b10100000_0111_011: DATA = 1'b0;
            15'b10100000_0111_100: DATA = 1'b0;
            15'b10100000_0111_101: DATA = 1'b0;
            15'b10100000_0111_110: DATA = 1'b0;
            15'b10100000_0111_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 2 Row 8
            15'b10100000_1000_000: DATA = 1'b0;
            15'b10100000_1000_001: DATA = 1'b0;
            15'b10100000_1000_010: DATA = 1'b0;
            15'b10100000_1000_011: DATA = 1'b0;
            15'b10100000_1000_100: DATA = 1'b0;
            15'b10100000_1000_101: DATA = 1'b0;
            15'b10100000_1000_110: DATA = 1'b0;
            15'b10100000_1000_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 2 Row 9
            15'b10100000_1001_000: DATA = 1'b0;
            15'b10100000_1001_001: DATA = 1'b0;
            15'b10100000_1001_010: DATA = 1'b0;
            15'b10100000_1001_011: DATA = 1'b0;
            15'b10100000_1001_100: DATA = 1'b0;
            15'b10100000_1001_101: DATA = 1'b0;
            15'b10100000_1001_110: DATA = 1'b0;
            15'b10100000_1001_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 2 Row 10
            15'b10100000_1010_000: DATA = 1'b0;
            15'b10100000_1010_001: DATA = 1'b0;
            15'b10100000_1010_010: DATA = 1'b0;
            15'b10100000_1010_011: DATA = 1'b0;
            15'b10100000_1010_100: DATA = 1'b0;
            15'b10100000_1010_101: DATA = 1'b0;
            15'b10100000_1010_110: DATA = 1'b0;
            15'b10100000_1010_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 2 Row 11
            15'b10100000_1011_000: DATA = 1'b0;
            15'b10100000_1011_001: DATA = 1'b0;
            15'b10100000_1011_010: DATA = 1'b0;
            15'b10100000_1011_011: DATA = 1'b0;
            15'b10100000_1011_100: DATA = 1'b0;
            15'b10100000_1011_101: DATA = 1'b0;
            15'b10100000_1011_110: DATA = 1'b0;
            15'b10100000_1011_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 2 Row 12
            15'b10100000_1100_000: DATA = 1'b0;
            15'b10100000_1100_001: DATA = 1'b0;
            15'b10100000_1100_010: DATA = 1'b0;
            15'b10100000_1100_011: DATA = 1'b0;
            15'b10100000_1100_100: DATA = 1'b0;
            15'b10100000_1100_101: DATA = 1'b0;
            15'b10100000_1100_110: DATA = 1'b0;
            15'b10100000_1100_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 2 Row 13
            15'b10100000_1101_000: DATA = 1'b0;
            15'b10100000_1101_001: DATA = 1'b0;
            15'b10100000_1101_010: DATA = 1'b0;
            15'b10100000_1101_011: DATA = 1'b0;
            15'b10100000_1101_100: DATA = 1'b0;
            15'b10100000_1101_101: DATA = 1'b0;
            15'b10100000_1101_110: DATA = 1'b0;
            15'b10100000_1101_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 2 Row 14
            15'b10100000_1110_000: DATA = 1'b0;
            15'b10100000_1110_001: DATA = 1'b0;
            15'b10100000_1110_010: DATA = 1'b0;
            15'b10100000_1110_011: DATA = 1'b0;
            15'b10100000_1110_100: DATA = 1'b0;
            15'b10100000_1110_101: DATA = 1'b0;
            15'b10100000_1110_110: DATA = 1'b0;
            15'b10100000_1110_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 2 Row 15
            15'b10100000_1111_000: DATA = 1'b0;
            15'b10100000_1111_001: DATA = 1'b0;
            15'b10100000_1111_010: DATA = 1'b0;
            15'b10100000_1111_011: DATA = 1'b0;
            15'b10100000_1111_100: DATA = 1'b0;
            15'b10100000_1111_101: DATA = 1'b0;
            15'b10100000_1111_110: DATA = 1'b0;
            15'b10100000_1111_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 3 Row 0
            15'b10100001_0000_000: DATA = 1'b0;
            15'b10100001_0000_001: DATA = 1'b0;
            15'b10100001_0000_010: DATA = 1'b0;
            15'b10100001_0000_011: DATA = 1'b0;
            15'b10100001_0000_100: DATA = 1'b0;
            15'b10100001_0000_101: DATA = 1'b0;
            15'b10100001_0000_110: DATA = 1'b0;
            15'b10100001_0000_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 3 Row 1
            15'b10100001_0001_000: DATA = 1'b0;
            15'b10100001_0001_001: DATA = 1'b0;
            15'b10100001_0001_010: DATA = 1'b0;
            15'b10100001_0001_011: DATA = 1'b0;
            15'b10100001_0001_100: DATA = 1'b0;
            15'b10100001_0001_101: DATA = 1'b0;
            15'b10100001_0001_110: DATA = 1'b0;
            15'b10100001_0001_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 3 Row 2
            15'b10100001_0010_000: DATA = 1'b0;
            15'b10100001_0010_001: DATA = 1'b0;
            15'b10100001_0010_010: DATA = 1'b0;
            15'b10100001_0010_011: DATA = 1'b0;
            15'b10100001_0010_100: DATA = 1'b0;
            15'b10100001_0010_101: DATA = 1'b0;
            15'b10100001_0010_110: DATA = 1'b0;
            15'b10100001_0010_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 3 Row 3
            15'b10100001_0011_000: DATA = 1'b0;
            15'b10100001_0011_001: DATA = 1'b0;
            15'b10100001_0011_010: DATA = 1'b0;
            15'b10100001_0011_011: DATA = 1'b0;
            15'b10100001_0011_100: DATA = 1'b0;
            15'b10100001_0011_101: DATA = 1'b0;
            15'b10100001_0011_110: DATA = 1'b0;
            15'b10100001_0011_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 3 Row 4
            15'b10100001_0100_000: DATA = 1'b0;
            15'b10100001_0100_001: DATA = 1'b0;
            15'b10100001_0100_010: DATA = 1'b0;
            15'b10100001_0100_011: DATA = 1'b0;
            15'b10100001_0100_100: DATA = 1'b0;
            15'b10100001_0100_101: DATA = 1'b0;
            15'b10100001_0100_110: DATA = 1'b0;
            15'b10100001_0100_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 3 Row 5
            15'b10100001_0101_000: DATA = 1'b0;
            15'b10100001_0101_001: DATA = 1'b0;
            15'b10100001_0101_010: DATA = 1'b0;
            15'b10100001_0101_011: DATA = 1'b0;
            15'b10100001_0101_100: DATA = 1'b0;
            15'b10100001_0101_101: DATA = 1'b0;
            15'b10100001_0101_110: DATA = 1'b0;
            15'b10100001_0101_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 3 Row 6
            15'b10100001_0110_000: DATA = 1'b0;
            15'b10100001_0110_001: DATA = 1'b0;
            15'b10100001_0110_010: DATA = 1'b0;
            15'b10100001_0110_011: DATA = 1'b0;
            15'b10100001_0110_100: DATA = 1'b0;
            15'b10100001_0110_101: DATA = 1'b0;
            15'b10100001_0110_110: DATA = 1'b0;
            15'b10100001_0110_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 3 Row 7
            15'b10100001_0111_000: DATA = 1'b0;
            15'b10100001_0111_001: DATA = 1'b0;
            15'b10100001_0111_010: DATA = 1'b0;
            15'b10100001_0111_011: DATA = 1'b0;
            15'b10100001_0111_100: DATA = 1'b0;
            15'b10100001_0111_101: DATA = 1'b0;
            15'b10100001_0111_110: DATA = 1'b0;
            15'b10100001_0111_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 3 Row 8
            15'b10100001_1000_000: DATA = 1'b0;
            15'b10100001_1000_001: DATA = 1'b0;
            15'b10100001_1000_010: DATA = 1'b0;
            15'b10100001_1000_011: DATA = 1'b0;
            15'b10100001_1000_100: DATA = 1'b0;
            15'b10100001_1000_101: DATA = 1'b0;
            15'b10100001_1000_110: DATA = 1'b0;
            15'b10100001_1000_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 3 Row 9
            15'b10100001_1001_000: DATA = 1'b0;
            15'b10100001_1001_001: DATA = 1'b0;
            15'b10100001_1001_010: DATA = 1'b0;
            15'b10100001_1001_011: DATA = 1'b0;
            15'b10100001_1001_100: DATA = 1'b0;
            15'b10100001_1001_101: DATA = 1'b0;
            15'b10100001_1001_110: DATA = 1'b0;
            15'b10100001_1001_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 3 Row 10
            15'b10100001_1010_000: DATA = 1'b0;
            15'b10100001_1010_001: DATA = 1'b0;
            15'b10100001_1010_010: DATA = 1'b0;
            15'b10100001_1010_011: DATA = 1'b0;
            15'b10100001_1010_100: DATA = 1'b0;
            15'b10100001_1010_101: DATA = 1'b0;
            15'b10100001_1010_110: DATA = 1'b0;
            15'b10100001_1010_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 3 Row 11
            15'b10100001_1011_000: DATA = 1'b0;
            15'b10100001_1011_001: DATA = 1'b0;
            15'b10100001_1011_010: DATA = 1'b0;
            15'b10100001_1011_011: DATA = 1'b0;
            15'b10100001_1011_100: DATA = 1'b0;
            15'b10100001_1011_101: DATA = 1'b0;
            15'b10100001_1011_110: DATA = 1'b0;
            15'b10100001_1011_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 3 Row 12
            15'b10100001_1100_000: DATA = 1'b0;
            15'b10100001_1100_001: DATA = 1'b0;
            15'b10100001_1100_010: DATA = 1'b0;
            15'b10100001_1100_011: DATA = 1'b0;
            15'b10100001_1100_100: DATA = 1'b0;
            15'b10100001_1100_101: DATA = 1'b0;
            15'b10100001_1100_110: DATA = 1'b0;
            15'b10100001_1100_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 3 Row 13
            15'b10100001_1101_000: DATA = 1'b0;
            15'b10100001_1101_001: DATA = 1'b0;
            15'b10100001_1101_010: DATA = 1'b0;
            15'b10100001_1101_011: DATA = 1'b0;
            15'b10100001_1101_100: DATA = 1'b0;
            15'b10100001_1101_101: DATA = 1'b0;
            15'b10100001_1101_110: DATA = 1'b0;
            15'b10100001_1101_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 3 Row 14
            15'b10100001_1110_000: DATA = 1'b0;
            15'b10100001_1110_001: DATA = 1'b0;
            15'b10100001_1110_010: DATA = 1'b0;
            15'b10100001_1110_011: DATA = 1'b0;
            15'b10100001_1110_100: DATA = 1'b0;
            15'b10100001_1110_101: DATA = 1'b0;
            15'b10100001_1110_110: DATA = 1'b0;
            15'b10100001_1110_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 3 Row 15
            15'b10100001_1111_000: DATA = 1'b0;
            15'b10100001_1111_001: DATA = 1'b0;
            15'b10100001_1111_010: DATA = 1'b0;
            15'b10100001_1111_011: DATA = 1'b0;
            15'b10100001_1111_100: DATA = 1'b0;
            15'b10100001_1111_101: DATA = 1'b0;
            15'b10100001_1111_110: DATA = 1'b0;
            15'b10100001_1111_111: DATA = 1'b0;
            // SQUARE- ROW 0 COL 4 Row 0
            15'b10100010_0000_000: DATA = 1'b0;
            15'b10100010_0000_001: DATA = 1'b0;
            15'b10100010_0000_010: DATA = 1'b0;
            15'b10100010_0000_011: DATA = 1'b0;
            15'b10100010_0000_100: DATA = 1'b0;
            15'b10100010_0000_101: DATA = 1'b0;
            15'b10100010_0000_110: DATA = 1'b0;
            15'b10100010_0000_111: DATA = 1'b1;
            // SQUARE- ROW 0 COL 4 Row 1
            15'b10100010_0001_000: DATA = 1'b0;
            15'b10100010_0001_001: DATA = 1'b0;
            15'b10100010_0001_010: DATA = 1'b0;
            15'b10100010_0001_011: DATA = 1'b0;
            15'b10100010_0001_100: DATA = 1'b0;
            15'b10100010_0001_101: DATA = 1'b0;
            15'b10100010_0001_110: DATA = 1'b0;
            15'b10100010_0001_111: DATA = 1'b1;
            // SQUARE- ROW 0 COL 4 Row 2
            15'b10100010_0010_000: DATA = 1'b0;
            15'b10100010_0010_001: DATA = 1'b0;
            15'b10100010_0010_010: DATA = 1'b0;
            15'b10100010_0010_011: DATA = 1'b0;
            15'b10100010_0010_100: DATA = 1'b0;
            15'b10100010_0010_101: DATA = 1'b0;
            15'b10100010_0010_110: DATA = 1'b0;
            15'b10100010_0010_111: DATA = 1'b1;
            // SQUARE- ROW 0 COL 4 Row 3
            15'b10100010_0011_000: DATA = 1'b0;
            15'b10100010_0011_001: DATA = 1'b0;
            15'b10100010_0011_010: DATA = 1'b0;
            15'b10100010_0011_011: DATA = 1'b0;
            15'b10100010_0011_100: DATA = 1'b0;
            15'b10100010_0011_101: DATA = 1'b0;
            15'b10100010_0011_110: DATA = 1'b0;
            15'b10100010_0011_111: DATA = 1'b1;
            // SQUARE- ROW 0 COL 4 Row 4
            15'b10100010_0100_000: DATA = 1'b0;
            15'b10100010_0100_001: DATA = 1'b0;
            15'b10100010_0100_010: DATA = 1'b0;
            15'b10100010_0100_011: DATA = 1'b0;
            15'b10100010_0100_100: DATA = 1'b0;
            15'b10100010_0100_101: DATA = 1'b0;
            15'b10100010_0100_110: DATA = 1'b0;
            15'b10100010_0100_111: DATA = 1'b1;
            // SQUARE- ROW 0 COL 4 Row 5
            15'b10100010_0101_000: DATA = 1'b0;
            15'b10100010_0101_001: DATA = 1'b0;
            15'b10100010_0101_010: DATA = 1'b0;
            15'b10100010_0101_011: DATA = 1'b0;
            15'b10100010_0101_100: DATA = 1'b0;
            15'b10100010_0101_101: DATA = 1'b0;
            15'b10100010_0101_110: DATA = 1'b0;
            15'b10100010_0101_111: DATA = 1'b1;
            // SQUARE- ROW 0 COL 4 Row 6
            15'b10100010_0110_000: DATA = 1'b0;
            15'b10100010_0110_001: DATA = 1'b0;
            15'b10100010_0110_010: DATA = 1'b0;
            15'b10100010_0110_011: DATA = 1'b0;
            15'b10100010_0110_100: DATA = 1'b0;
            15'b10100010_0110_101: DATA = 1'b0;
            15'b10100010_0110_110: DATA = 1'b0;
            15'b10100010_0110_111: DATA = 1'b1;
            // SQUARE- ROW 0 COL 4 Row 7
            15'b10100010_0111_000: DATA = 1'b0;
            15'b10100010_0111_001: DATA = 1'b0;
            15'b10100010_0111_010: DATA = 1'b0;
            15'b10100010_0111_011: DATA = 1'b0;
            15'b10100010_0111_100: DATA = 1'b0;
            15'b10100010_0111_101: DATA = 1'b0;
            15'b10100010_0111_110: DATA = 1'b0;
            15'b10100010_0111_111: DATA = 1'b1;
            // SQUARE- ROW 0 COL 4 Row 8
            15'b10100010_1000_000: DATA = 1'b0;
            15'b10100010_1000_001: DATA = 1'b0;
            15'b10100010_1000_010: DATA = 1'b0;
            15'b10100010_1000_011: DATA = 1'b0;
            15'b10100010_1000_100: DATA = 1'b0;
            15'b10100010_1000_101: DATA = 1'b0;
            15'b10100010_1000_110: DATA = 1'b0;
            15'b10100010_1000_111: DATA = 1'b1;
            // SQUARE- ROW 0 COL 4 Row 9
            15'b10100010_1001_000: DATA = 1'b0;
            15'b10100010_1001_001: DATA = 1'b0;
            15'b10100010_1001_010: DATA = 1'b0;
            15'b10100010_1001_011: DATA = 1'b0;
            15'b10100010_1001_100: DATA = 1'b0;
            15'b10100010_1001_101: DATA = 1'b0;
            15'b10100010_1001_110: DATA = 1'b0;
            15'b10100010_1001_111: DATA = 1'b1;
            // SQUARE- ROW 0 COL 4 Row 10
            15'b10100010_1010_000: DATA = 1'b0;
            15'b10100010_1010_001: DATA = 1'b0;
            15'b10100010_1010_010: DATA = 1'b0;
            15'b10100010_1010_011: DATA = 1'b0;
            15'b10100010_1010_100: DATA = 1'b0;
            15'b10100010_1010_101: DATA = 1'b0;
            15'b10100010_1010_110: DATA = 1'b0;
            15'b10100010_1010_111: DATA = 1'b1;
            // SQUARE- ROW 0 COL 4 Row 11
            15'b10100010_1011_000: DATA = 1'b0;
            15'b10100010_1011_001: DATA = 1'b0;
            15'b10100010_1011_010: DATA = 1'b0;
            15'b10100010_1011_011: DATA = 1'b0;
            15'b10100010_1011_100: DATA = 1'b0;
            15'b10100010_1011_101: DATA = 1'b0;
            15'b10100010_1011_110: DATA = 1'b0;
            15'b10100010_1011_111: DATA = 1'b1;
            // SQUARE- ROW 0 COL 4 Row 12
            15'b10100010_1100_000: DATA = 1'b0;
            15'b10100010_1100_001: DATA = 1'b0;
            15'b10100010_1100_010: DATA = 1'b0;
            15'b10100010_1100_011: DATA = 1'b0;
            15'b10100010_1100_100: DATA = 1'b0;
            15'b10100010_1100_101: DATA = 1'b0;
            15'b10100010_1100_110: DATA = 1'b0;
            15'b10100010_1100_111: DATA = 1'b1;
            // SQUARE- ROW 0 COL 4 Row 13
            15'b10100010_1101_000: DATA = 1'b0;
            15'b10100010_1101_001: DATA = 1'b0;
            15'b10100010_1101_010: DATA = 1'b0;
            15'b10100010_1101_011: DATA = 1'b0;
            15'b10100010_1101_100: DATA = 1'b0;
            15'b10100010_1101_101: DATA = 1'b0;
            15'b10100010_1101_110: DATA = 1'b0;
            15'b10100010_1101_111: DATA = 1'b1;
            // SQUARE- ROW 0 COL 4 Row 14
            15'b10100010_1110_000: DATA = 1'b0;
            15'b10100010_1110_001: DATA = 1'b0;
            15'b10100010_1110_010: DATA = 1'b0;
            15'b10100010_1110_011: DATA = 1'b0;
            15'b10100010_1110_100: DATA = 1'b0;
            15'b10100010_1110_101: DATA = 1'b0;
            15'b10100010_1110_110: DATA = 1'b0;
            15'b10100010_1110_111: DATA = 1'b1;
            // SQUARE- ROW 0 COL 4 Row 15
            15'b10100010_1111_000: DATA = 1'b0;
            15'b10100010_1111_001: DATA = 1'b0;
            15'b10100010_1111_010: DATA = 1'b0;
            15'b10100010_1111_011: DATA = 1'b0;
            15'b10100010_1111_100: DATA = 1'b0;
            15'b10100010_1111_101: DATA = 1'b0;
            15'b10100010_1111_110: DATA = 1'b0;
            15'b10100010_1111_111: DATA = 1'b1;
            // SQUARE- ROW 1 COL 0 Row 0
            15'b10100011_0000_000: DATA = 1'b1;
            15'b10100011_0000_001: DATA = 1'b0;
            15'b10100011_0000_010: DATA = 1'b0;
            15'b10100011_0000_011: DATA = 1'b0;
            15'b10100011_0000_100: DATA = 1'b0;
            15'b10100011_0000_101: DATA = 1'b0;
            15'b10100011_0000_110: DATA = 1'b0;
            15'b10100011_0000_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 0 Row 1
            15'b10100011_0001_000: DATA = 1'b1;
            15'b10100011_0001_001: DATA = 1'b0;
            15'b10100011_0001_010: DATA = 1'b0;
            15'b10100011_0001_011: DATA = 1'b0;
            15'b10100011_0001_100: DATA = 1'b0;
            15'b10100011_0001_101: DATA = 1'b0;
            15'b10100011_0001_110: DATA = 1'b0;
            15'b10100011_0001_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 0 Row 2
            15'b10100011_0010_000: DATA = 1'b1;
            15'b10100011_0010_001: DATA = 1'b0;
            15'b10100011_0010_010: DATA = 1'b0;
            15'b10100011_0010_011: DATA = 1'b0;
            15'b10100011_0010_100: DATA = 1'b0;
            15'b10100011_0010_101: DATA = 1'b0;
            15'b10100011_0010_110: DATA = 1'b0;
            15'b10100011_0010_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 0 Row 3
            15'b10100011_0011_000: DATA = 1'b1;
            15'b10100011_0011_001: DATA = 1'b0;
            15'b10100011_0011_010: DATA = 1'b0;
            15'b10100011_0011_011: DATA = 1'b0;
            15'b10100011_0011_100: DATA = 1'b0;
            15'b10100011_0011_101: DATA = 1'b0;
            15'b10100011_0011_110: DATA = 1'b0;
            15'b10100011_0011_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 0 Row 4
            15'b10100011_0100_000: DATA = 1'b1;
            15'b10100011_0100_001: DATA = 1'b0;
            15'b10100011_0100_010: DATA = 1'b0;
            15'b10100011_0100_011: DATA = 1'b0;
            15'b10100011_0100_100: DATA = 1'b0;
            15'b10100011_0100_101: DATA = 1'b0;
            15'b10100011_0100_110: DATA = 1'b0;
            15'b10100011_0100_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 0 Row 5
            15'b10100011_0101_000: DATA = 1'b1;
            15'b10100011_0101_001: DATA = 1'b0;
            15'b10100011_0101_010: DATA = 1'b0;
            15'b10100011_0101_011: DATA = 1'b0;
            15'b10100011_0101_100: DATA = 1'b0;
            15'b10100011_0101_101: DATA = 1'b0;
            15'b10100011_0101_110: DATA = 1'b0;
            15'b10100011_0101_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 0 Row 6
            15'b10100011_0110_000: DATA = 1'b1;
            15'b10100011_0110_001: DATA = 1'b0;
            15'b10100011_0110_010: DATA = 1'b0;
            15'b10100011_0110_011: DATA = 1'b0;
            15'b10100011_0110_100: DATA = 1'b0;
            15'b10100011_0110_101: DATA = 1'b0;
            15'b10100011_0110_110: DATA = 1'b0;
            15'b10100011_0110_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 0 Row 7
            15'b10100011_0111_000: DATA = 1'b1;
            15'b10100011_0111_001: DATA = 1'b0;
            15'b10100011_0111_010: DATA = 1'b0;
            15'b10100011_0111_011: DATA = 1'b0;
            15'b10100011_0111_100: DATA = 1'b0;
            15'b10100011_0111_101: DATA = 1'b0;
            15'b10100011_0111_110: DATA = 1'b0;
            15'b10100011_0111_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 0 Row 8
            15'b10100011_1000_000: DATA = 1'b1;
            15'b10100011_1000_001: DATA = 1'b0;
            15'b10100011_1000_010: DATA = 1'b0;
            15'b10100011_1000_011: DATA = 1'b0;
            15'b10100011_1000_100: DATA = 1'b0;
            15'b10100011_1000_101: DATA = 1'b0;
            15'b10100011_1000_110: DATA = 1'b0;
            15'b10100011_1000_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 0 Row 9
            15'b10100011_1001_000: DATA = 1'b1;
            15'b10100011_1001_001: DATA = 1'b0;
            15'b10100011_1001_010: DATA = 1'b0;
            15'b10100011_1001_011: DATA = 1'b0;
            15'b10100011_1001_100: DATA = 1'b0;
            15'b10100011_1001_101: DATA = 1'b0;
            15'b10100011_1001_110: DATA = 1'b0;
            15'b10100011_1001_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 0 Row 10
            15'b10100011_1010_000: DATA = 1'b1;
            15'b10100011_1010_001: DATA = 1'b0;
            15'b10100011_1010_010: DATA = 1'b0;
            15'b10100011_1010_011: DATA = 1'b0;
            15'b10100011_1010_100: DATA = 1'b0;
            15'b10100011_1010_101: DATA = 1'b0;
            15'b10100011_1010_110: DATA = 1'b0;
            15'b10100011_1010_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 0 Row 11
            15'b10100011_1011_000: DATA = 1'b1;
            15'b10100011_1011_001: DATA = 1'b0;
            15'b10100011_1011_010: DATA = 1'b0;
            15'b10100011_1011_011: DATA = 1'b0;
            15'b10100011_1011_100: DATA = 1'b0;
            15'b10100011_1011_101: DATA = 1'b0;
            15'b10100011_1011_110: DATA = 1'b0;
            15'b10100011_1011_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 0 Row 12
            15'b10100011_1100_000: DATA = 1'b1;
            15'b10100011_1100_001: DATA = 1'b0;
            15'b10100011_1100_010: DATA = 1'b0;
            15'b10100011_1100_011: DATA = 1'b0;
            15'b10100011_1100_100: DATA = 1'b0;
            15'b10100011_1100_101: DATA = 1'b0;
            15'b10100011_1100_110: DATA = 1'b0;
            15'b10100011_1100_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 0 Row 13
            15'b10100011_1101_000: DATA = 1'b1;
            15'b10100011_1101_001: DATA = 1'b0;
            15'b10100011_1101_010: DATA = 1'b0;
            15'b10100011_1101_011: DATA = 1'b0;
            15'b10100011_1101_100: DATA = 1'b0;
            15'b10100011_1101_101: DATA = 1'b0;
            15'b10100011_1101_110: DATA = 1'b0;
            15'b10100011_1101_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 0 Row 14
            15'b10100011_1110_000: DATA = 1'b1;
            15'b10100011_1110_001: DATA = 1'b0;
            15'b10100011_1110_010: DATA = 1'b0;
            15'b10100011_1110_011: DATA = 1'b0;
            15'b10100011_1110_100: DATA = 1'b0;
            15'b10100011_1110_101: DATA = 1'b0;
            15'b10100011_1110_110: DATA = 1'b0;
            15'b10100011_1110_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 0 Row 15
            15'b10100011_1111_000: DATA = 1'b1;
            15'b10100011_1111_001: DATA = 1'b1;
            15'b10100011_1111_010: DATA = 1'b1;
            15'b10100011_1111_011: DATA = 1'b1;
            15'b10100011_1111_100: DATA = 1'b1;
            15'b10100011_1111_101: DATA = 1'b1;
            15'b10100011_1111_110: DATA = 1'b1;
            15'b10100011_1111_111: DATA = 1'b1;
            // SQUARE- ROW 1 COL 1 Row 0
            15'b10100100_0000_000: DATA = 1'b0;
            15'b10100100_0000_001: DATA = 1'b0;
            15'b10100100_0000_010: DATA = 1'b0;
            15'b10100100_0000_011: DATA = 1'b0;
            15'b10100100_0000_100: DATA = 1'b0;
            15'b10100100_0000_101: DATA = 1'b0;
            15'b10100100_0000_110: DATA = 1'b0;
            15'b10100100_0000_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 1 Row 1
            15'b10100100_0001_000: DATA = 1'b0;
            15'b10100100_0001_001: DATA = 1'b0;
            15'b10100100_0001_010: DATA = 1'b0;
            15'b10100100_0001_011: DATA = 1'b0;
            15'b10100100_0001_100: DATA = 1'b0;
            15'b10100100_0001_101: DATA = 1'b0;
            15'b10100100_0001_110: DATA = 1'b0;
            15'b10100100_0001_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 1 Row 2
            15'b10100100_0010_000: DATA = 1'b0;
            15'b10100100_0010_001: DATA = 1'b0;
            15'b10100100_0010_010: DATA = 1'b0;
            15'b10100100_0010_011: DATA = 1'b0;
            15'b10100100_0010_100: DATA = 1'b0;
            15'b10100100_0010_101: DATA = 1'b0;
            15'b10100100_0010_110: DATA = 1'b0;
            15'b10100100_0010_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 1 Row 3
            15'b10100100_0011_000: DATA = 1'b0;
            15'b10100100_0011_001: DATA = 1'b0;
            15'b10100100_0011_010: DATA = 1'b0;
            15'b10100100_0011_011: DATA = 1'b0;
            15'b10100100_0011_100: DATA = 1'b0;
            15'b10100100_0011_101: DATA = 1'b0;
            15'b10100100_0011_110: DATA = 1'b0;
            15'b10100100_0011_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 1 Row 4
            15'b10100100_0100_000: DATA = 1'b0;
            15'b10100100_0100_001: DATA = 1'b0;
            15'b10100100_0100_010: DATA = 1'b0;
            15'b10100100_0100_011: DATA = 1'b0;
            15'b10100100_0100_100: DATA = 1'b0;
            15'b10100100_0100_101: DATA = 1'b0;
            15'b10100100_0100_110: DATA = 1'b0;
            15'b10100100_0100_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 1 Row 5
            15'b10100100_0101_000: DATA = 1'b0;
            15'b10100100_0101_001: DATA = 1'b0;
            15'b10100100_0101_010: DATA = 1'b0;
            15'b10100100_0101_011: DATA = 1'b0;
            15'b10100100_0101_100: DATA = 1'b0;
            15'b10100100_0101_101: DATA = 1'b0;
            15'b10100100_0101_110: DATA = 1'b0;
            15'b10100100_0101_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 1 Row 6
            15'b10100100_0110_000: DATA = 1'b0;
            15'b10100100_0110_001: DATA = 1'b0;
            15'b10100100_0110_010: DATA = 1'b0;
            15'b10100100_0110_011: DATA = 1'b0;
            15'b10100100_0110_100: DATA = 1'b0;
            15'b10100100_0110_101: DATA = 1'b0;
            15'b10100100_0110_110: DATA = 1'b0;
            15'b10100100_0110_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 1 Row 7
            15'b10100100_0111_000: DATA = 1'b0;
            15'b10100100_0111_001: DATA = 1'b0;
            15'b10100100_0111_010: DATA = 1'b0;
            15'b10100100_0111_011: DATA = 1'b0;
            15'b10100100_0111_100: DATA = 1'b0;
            15'b10100100_0111_101: DATA = 1'b0;
            15'b10100100_0111_110: DATA = 1'b0;
            15'b10100100_0111_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 1 Row 8
            15'b10100100_1000_000: DATA = 1'b0;
            15'b10100100_1000_001: DATA = 1'b0;
            15'b10100100_1000_010: DATA = 1'b0;
            15'b10100100_1000_011: DATA = 1'b0;
            15'b10100100_1000_100: DATA = 1'b0;
            15'b10100100_1000_101: DATA = 1'b0;
            15'b10100100_1000_110: DATA = 1'b0;
            15'b10100100_1000_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 1 Row 9
            15'b10100100_1001_000: DATA = 1'b0;
            15'b10100100_1001_001: DATA = 1'b0;
            15'b10100100_1001_010: DATA = 1'b0;
            15'b10100100_1001_011: DATA = 1'b0;
            15'b10100100_1001_100: DATA = 1'b0;
            15'b10100100_1001_101: DATA = 1'b0;
            15'b10100100_1001_110: DATA = 1'b0;
            15'b10100100_1001_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 1 Row 10
            15'b10100100_1010_000: DATA = 1'b0;
            15'b10100100_1010_001: DATA = 1'b0;
            15'b10100100_1010_010: DATA = 1'b0;
            15'b10100100_1010_011: DATA = 1'b0;
            15'b10100100_1010_100: DATA = 1'b0;
            15'b10100100_1010_101: DATA = 1'b0;
            15'b10100100_1010_110: DATA = 1'b0;
            15'b10100100_1010_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 1 Row 11
            15'b10100100_1011_000: DATA = 1'b0;
            15'b10100100_1011_001: DATA = 1'b0;
            15'b10100100_1011_010: DATA = 1'b0;
            15'b10100100_1011_011: DATA = 1'b0;
            15'b10100100_1011_100: DATA = 1'b0;
            15'b10100100_1011_101: DATA = 1'b0;
            15'b10100100_1011_110: DATA = 1'b0;
            15'b10100100_1011_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 1 Row 12
            15'b10100100_1100_000: DATA = 1'b0;
            15'b10100100_1100_001: DATA = 1'b0;
            15'b10100100_1100_010: DATA = 1'b0;
            15'b10100100_1100_011: DATA = 1'b0;
            15'b10100100_1100_100: DATA = 1'b0;
            15'b10100100_1100_101: DATA = 1'b0;
            15'b10100100_1100_110: DATA = 1'b0;
            15'b10100100_1100_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 1 Row 13
            15'b10100100_1101_000: DATA = 1'b0;
            15'b10100100_1101_001: DATA = 1'b0;
            15'b10100100_1101_010: DATA = 1'b0;
            15'b10100100_1101_011: DATA = 1'b0;
            15'b10100100_1101_100: DATA = 1'b0;
            15'b10100100_1101_101: DATA = 1'b0;
            15'b10100100_1101_110: DATA = 1'b0;
            15'b10100100_1101_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 1 Row 14
            15'b10100100_1110_000: DATA = 1'b0;
            15'b10100100_1110_001: DATA = 1'b0;
            15'b10100100_1110_010: DATA = 1'b0;
            15'b10100100_1110_011: DATA = 1'b0;
            15'b10100100_1110_100: DATA = 1'b0;
            15'b10100100_1110_101: DATA = 1'b0;
            15'b10100100_1110_110: DATA = 1'b0;
            15'b10100100_1110_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 1 Row 15
            15'b10100100_1111_000: DATA = 1'b1;
            15'b10100100_1111_001: DATA = 1'b1;
            15'b10100100_1111_010: DATA = 1'b1;
            15'b10100100_1111_011: DATA = 1'b1;
            15'b10100100_1111_100: DATA = 1'b1;
            15'b10100100_1111_101: DATA = 1'b1;
            15'b10100100_1111_110: DATA = 1'b1;
            15'b10100100_1111_111: DATA = 1'b1;
            // SQUARE- ROW 1 COL 2 Row 0
            15'b10100101_0000_000: DATA = 1'b0;
            15'b10100101_0000_001: DATA = 1'b0;
            15'b10100101_0000_010: DATA = 1'b0;
            15'b10100101_0000_011: DATA = 1'b0;
            15'b10100101_0000_100: DATA = 1'b0;
            15'b10100101_0000_101: DATA = 1'b0;
            15'b10100101_0000_110: DATA = 1'b0;
            15'b10100101_0000_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 2 Row 1
            15'b10100101_0001_000: DATA = 1'b0;
            15'b10100101_0001_001: DATA = 1'b0;
            15'b10100101_0001_010: DATA = 1'b0;
            15'b10100101_0001_011: DATA = 1'b0;
            15'b10100101_0001_100: DATA = 1'b0;
            15'b10100101_0001_101: DATA = 1'b0;
            15'b10100101_0001_110: DATA = 1'b0;
            15'b10100101_0001_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 2 Row 2
            15'b10100101_0010_000: DATA = 1'b0;
            15'b10100101_0010_001: DATA = 1'b0;
            15'b10100101_0010_010: DATA = 1'b0;
            15'b10100101_0010_011: DATA = 1'b0;
            15'b10100101_0010_100: DATA = 1'b0;
            15'b10100101_0010_101: DATA = 1'b0;
            15'b10100101_0010_110: DATA = 1'b0;
            15'b10100101_0010_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 2 Row 3
            15'b10100101_0011_000: DATA = 1'b0;
            15'b10100101_0011_001: DATA = 1'b0;
            15'b10100101_0011_010: DATA = 1'b0;
            15'b10100101_0011_011: DATA = 1'b0;
            15'b10100101_0011_100: DATA = 1'b0;
            15'b10100101_0011_101: DATA = 1'b0;
            15'b10100101_0011_110: DATA = 1'b0;
            15'b10100101_0011_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 2 Row 4
            15'b10100101_0100_000: DATA = 1'b0;
            15'b10100101_0100_001: DATA = 1'b0;
            15'b10100101_0100_010: DATA = 1'b0;
            15'b10100101_0100_011: DATA = 1'b0;
            15'b10100101_0100_100: DATA = 1'b0;
            15'b10100101_0100_101: DATA = 1'b0;
            15'b10100101_0100_110: DATA = 1'b0;
            15'b10100101_0100_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 2 Row 5
            15'b10100101_0101_000: DATA = 1'b0;
            15'b10100101_0101_001: DATA = 1'b0;
            15'b10100101_0101_010: DATA = 1'b0;
            15'b10100101_0101_011: DATA = 1'b0;
            15'b10100101_0101_100: DATA = 1'b0;
            15'b10100101_0101_101: DATA = 1'b0;
            15'b10100101_0101_110: DATA = 1'b0;
            15'b10100101_0101_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 2 Row 6
            15'b10100101_0110_000: DATA = 1'b0;
            15'b10100101_0110_001: DATA = 1'b0;
            15'b10100101_0110_010: DATA = 1'b0;
            15'b10100101_0110_011: DATA = 1'b0;
            15'b10100101_0110_100: DATA = 1'b0;
            15'b10100101_0110_101: DATA = 1'b0;
            15'b10100101_0110_110: DATA = 1'b0;
            15'b10100101_0110_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 2 Row 7
            15'b10100101_0111_000: DATA = 1'b0;
            15'b10100101_0111_001: DATA = 1'b0;
            15'b10100101_0111_010: DATA = 1'b0;
            15'b10100101_0111_011: DATA = 1'b0;
            15'b10100101_0111_100: DATA = 1'b0;
            15'b10100101_0111_101: DATA = 1'b0;
            15'b10100101_0111_110: DATA = 1'b0;
            15'b10100101_0111_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 2 Row 8
            15'b10100101_1000_000: DATA = 1'b0;
            15'b10100101_1000_001: DATA = 1'b0;
            15'b10100101_1000_010: DATA = 1'b0;
            15'b10100101_1000_011: DATA = 1'b0;
            15'b10100101_1000_100: DATA = 1'b0;
            15'b10100101_1000_101: DATA = 1'b0;
            15'b10100101_1000_110: DATA = 1'b0;
            15'b10100101_1000_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 2 Row 9
            15'b10100101_1001_000: DATA = 1'b0;
            15'b10100101_1001_001: DATA = 1'b0;
            15'b10100101_1001_010: DATA = 1'b0;
            15'b10100101_1001_011: DATA = 1'b0;
            15'b10100101_1001_100: DATA = 1'b0;
            15'b10100101_1001_101: DATA = 1'b0;
            15'b10100101_1001_110: DATA = 1'b0;
            15'b10100101_1001_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 2 Row 10
            15'b10100101_1010_000: DATA = 1'b0;
            15'b10100101_1010_001: DATA = 1'b0;
            15'b10100101_1010_010: DATA = 1'b0;
            15'b10100101_1010_011: DATA = 1'b0;
            15'b10100101_1010_100: DATA = 1'b0;
            15'b10100101_1010_101: DATA = 1'b0;
            15'b10100101_1010_110: DATA = 1'b0;
            15'b10100101_1010_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 2 Row 11
            15'b10100101_1011_000: DATA = 1'b0;
            15'b10100101_1011_001: DATA = 1'b0;
            15'b10100101_1011_010: DATA = 1'b0;
            15'b10100101_1011_011: DATA = 1'b0;
            15'b10100101_1011_100: DATA = 1'b0;
            15'b10100101_1011_101: DATA = 1'b0;
            15'b10100101_1011_110: DATA = 1'b0;
            15'b10100101_1011_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 2 Row 12
            15'b10100101_1100_000: DATA = 1'b0;
            15'b10100101_1100_001: DATA = 1'b0;
            15'b10100101_1100_010: DATA = 1'b0;
            15'b10100101_1100_011: DATA = 1'b0;
            15'b10100101_1100_100: DATA = 1'b0;
            15'b10100101_1100_101: DATA = 1'b0;
            15'b10100101_1100_110: DATA = 1'b0;
            15'b10100101_1100_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 2 Row 13
            15'b10100101_1101_000: DATA = 1'b0;
            15'b10100101_1101_001: DATA = 1'b0;
            15'b10100101_1101_010: DATA = 1'b0;
            15'b10100101_1101_011: DATA = 1'b0;
            15'b10100101_1101_100: DATA = 1'b0;
            15'b10100101_1101_101: DATA = 1'b0;
            15'b10100101_1101_110: DATA = 1'b0;
            15'b10100101_1101_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 2 Row 14
            15'b10100101_1110_000: DATA = 1'b0;
            15'b10100101_1110_001: DATA = 1'b0;
            15'b10100101_1110_010: DATA = 1'b0;
            15'b10100101_1110_011: DATA = 1'b0;
            15'b10100101_1110_100: DATA = 1'b0;
            15'b10100101_1110_101: DATA = 1'b0;
            15'b10100101_1110_110: DATA = 1'b0;
            15'b10100101_1110_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 2 Row 15
            15'b10100101_1111_000: DATA = 1'b1;
            15'b10100101_1111_001: DATA = 1'b1;
            15'b10100101_1111_010: DATA = 1'b1;
            15'b10100101_1111_011: DATA = 1'b1;
            15'b10100101_1111_100: DATA = 1'b1;
            15'b10100101_1111_101: DATA = 1'b1;
            15'b10100101_1111_110: DATA = 1'b1;
            15'b10100101_1111_111: DATA = 1'b1;
            // SQUARE- ROW 1 COL 3 Row 0
            15'b10100110_0000_000: DATA = 1'b0;
            15'b10100110_0000_001: DATA = 1'b0;
            15'b10100110_0000_010: DATA = 1'b0;
            15'b10100110_0000_011: DATA = 1'b0;
            15'b10100110_0000_100: DATA = 1'b0;
            15'b10100110_0000_101: DATA = 1'b0;
            15'b10100110_0000_110: DATA = 1'b0;
            15'b10100110_0000_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 3 Row 1
            15'b10100110_0001_000: DATA = 1'b0;
            15'b10100110_0001_001: DATA = 1'b0;
            15'b10100110_0001_010: DATA = 1'b0;
            15'b10100110_0001_011: DATA = 1'b0;
            15'b10100110_0001_100: DATA = 1'b0;
            15'b10100110_0001_101: DATA = 1'b0;
            15'b10100110_0001_110: DATA = 1'b0;
            15'b10100110_0001_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 3 Row 2
            15'b10100110_0010_000: DATA = 1'b0;
            15'b10100110_0010_001: DATA = 1'b0;
            15'b10100110_0010_010: DATA = 1'b0;
            15'b10100110_0010_011: DATA = 1'b0;
            15'b10100110_0010_100: DATA = 1'b0;
            15'b10100110_0010_101: DATA = 1'b0;
            15'b10100110_0010_110: DATA = 1'b0;
            15'b10100110_0010_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 3 Row 3
            15'b10100110_0011_000: DATA = 1'b0;
            15'b10100110_0011_001: DATA = 1'b0;
            15'b10100110_0011_010: DATA = 1'b0;
            15'b10100110_0011_011: DATA = 1'b0;
            15'b10100110_0011_100: DATA = 1'b0;
            15'b10100110_0011_101: DATA = 1'b0;
            15'b10100110_0011_110: DATA = 1'b0;
            15'b10100110_0011_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 3 Row 4
            15'b10100110_0100_000: DATA = 1'b0;
            15'b10100110_0100_001: DATA = 1'b0;
            15'b10100110_0100_010: DATA = 1'b0;
            15'b10100110_0100_011: DATA = 1'b0;
            15'b10100110_0100_100: DATA = 1'b0;
            15'b10100110_0100_101: DATA = 1'b0;
            15'b10100110_0100_110: DATA = 1'b0;
            15'b10100110_0100_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 3 Row 5
            15'b10100110_0101_000: DATA = 1'b0;
            15'b10100110_0101_001: DATA = 1'b0;
            15'b10100110_0101_010: DATA = 1'b0;
            15'b10100110_0101_011: DATA = 1'b0;
            15'b10100110_0101_100: DATA = 1'b0;
            15'b10100110_0101_101: DATA = 1'b0;
            15'b10100110_0101_110: DATA = 1'b0;
            15'b10100110_0101_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 3 Row 6
            15'b10100110_0110_000: DATA = 1'b0;
            15'b10100110_0110_001: DATA = 1'b0;
            15'b10100110_0110_010: DATA = 1'b0;
            15'b10100110_0110_011: DATA = 1'b0;
            15'b10100110_0110_100: DATA = 1'b0;
            15'b10100110_0110_101: DATA = 1'b0;
            15'b10100110_0110_110: DATA = 1'b0;
            15'b10100110_0110_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 3 Row 7
            15'b10100110_0111_000: DATA = 1'b0;
            15'b10100110_0111_001: DATA = 1'b0;
            15'b10100110_0111_010: DATA = 1'b0;
            15'b10100110_0111_011: DATA = 1'b0;
            15'b10100110_0111_100: DATA = 1'b0;
            15'b10100110_0111_101: DATA = 1'b0;
            15'b10100110_0111_110: DATA = 1'b0;
            15'b10100110_0111_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 3 Row 8
            15'b10100110_1000_000: DATA = 1'b0;
            15'b10100110_1000_001: DATA = 1'b0;
            15'b10100110_1000_010: DATA = 1'b0;
            15'b10100110_1000_011: DATA = 1'b0;
            15'b10100110_1000_100: DATA = 1'b0;
            15'b10100110_1000_101: DATA = 1'b0;
            15'b10100110_1000_110: DATA = 1'b0;
            15'b10100110_1000_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 3 Row 9
            15'b10100110_1001_000: DATA = 1'b0;
            15'b10100110_1001_001: DATA = 1'b0;
            15'b10100110_1001_010: DATA = 1'b0;
            15'b10100110_1001_011: DATA = 1'b0;
            15'b10100110_1001_100: DATA = 1'b0;
            15'b10100110_1001_101: DATA = 1'b0;
            15'b10100110_1001_110: DATA = 1'b0;
            15'b10100110_1001_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 3 Row 10
            15'b10100110_1010_000: DATA = 1'b0;
            15'b10100110_1010_001: DATA = 1'b0;
            15'b10100110_1010_010: DATA = 1'b0;
            15'b10100110_1010_011: DATA = 1'b0;
            15'b10100110_1010_100: DATA = 1'b0;
            15'b10100110_1010_101: DATA = 1'b0;
            15'b10100110_1010_110: DATA = 1'b0;
            15'b10100110_1010_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 3 Row 11
            15'b10100110_1011_000: DATA = 1'b0;
            15'b10100110_1011_001: DATA = 1'b0;
            15'b10100110_1011_010: DATA = 1'b0;
            15'b10100110_1011_011: DATA = 1'b0;
            15'b10100110_1011_100: DATA = 1'b0;
            15'b10100110_1011_101: DATA = 1'b0;
            15'b10100110_1011_110: DATA = 1'b0;
            15'b10100110_1011_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 3 Row 12
            15'b10100110_1100_000: DATA = 1'b0;
            15'b10100110_1100_001: DATA = 1'b0;
            15'b10100110_1100_010: DATA = 1'b0;
            15'b10100110_1100_011: DATA = 1'b0;
            15'b10100110_1100_100: DATA = 1'b0;
            15'b10100110_1100_101: DATA = 1'b0;
            15'b10100110_1100_110: DATA = 1'b0;
            15'b10100110_1100_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 3 Row 13
            15'b10100110_1101_000: DATA = 1'b0;
            15'b10100110_1101_001: DATA = 1'b0;
            15'b10100110_1101_010: DATA = 1'b0;
            15'b10100110_1101_011: DATA = 1'b0;
            15'b10100110_1101_100: DATA = 1'b0;
            15'b10100110_1101_101: DATA = 1'b0;
            15'b10100110_1101_110: DATA = 1'b0;
            15'b10100110_1101_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 3 Row 14
            15'b10100110_1110_000: DATA = 1'b0;
            15'b10100110_1110_001: DATA = 1'b0;
            15'b10100110_1110_010: DATA = 1'b0;
            15'b10100110_1110_011: DATA = 1'b0;
            15'b10100110_1110_100: DATA = 1'b0;
            15'b10100110_1110_101: DATA = 1'b0;
            15'b10100110_1110_110: DATA = 1'b0;
            15'b10100110_1110_111: DATA = 1'b0;
            // SQUARE- ROW 1 COL 3 Row 15
            15'b10100110_1111_000: DATA = 1'b1;
            15'b10100110_1111_001: DATA = 1'b1;
            15'b10100110_1111_010: DATA = 1'b1;
            15'b10100110_1111_011: DATA = 1'b1;
            15'b10100110_1111_100: DATA = 1'b1;
            15'b10100110_1111_101: DATA = 1'b1;
            15'b10100110_1111_110: DATA = 1'b1;
            15'b10100110_1111_111: DATA = 1'b1;
            // SQUARE- ROW 1 COL 4 Row 0
            15'b10100111_0000_000: DATA = 1'b0;
            15'b10100111_0000_001: DATA = 1'b0;
            15'b10100111_0000_010: DATA = 1'b0;
            15'b10100111_0000_011: DATA = 1'b0;
            15'b10100111_0000_100: DATA = 1'b0;
            15'b10100111_0000_101: DATA = 1'b0;
            15'b10100111_0000_110: DATA = 1'b0;
            15'b10100111_0000_111: DATA = 1'b1;
            // SQUARE- ROW 1 COL 4 Row 1
            15'b10100111_0001_000: DATA = 1'b0;
            15'b10100111_0001_001: DATA = 1'b0;
            15'b10100111_0001_010: DATA = 1'b0;
            15'b10100111_0001_011: DATA = 1'b0;
            15'b10100111_0001_100: DATA = 1'b0;
            15'b10100111_0001_101: DATA = 1'b0;
            15'b10100111_0001_110: DATA = 1'b0;
            15'b10100111_0001_111: DATA = 1'b1;
            // SQUARE- ROW 1 COL 4 Row 2
            15'b10100111_0010_000: DATA = 1'b0;
            15'b10100111_0010_001: DATA = 1'b0;
            15'b10100111_0010_010: DATA = 1'b0;
            15'b10100111_0010_011: DATA = 1'b0;
            15'b10100111_0010_100: DATA = 1'b0;
            15'b10100111_0010_101: DATA = 1'b0;
            15'b10100111_0010_110: DATA = 1'b0;
            15'b10100111_0010_111: DATA = 1'b1;
            // SQUARE- ROW 1 COL 4 Row 3
            15'b10100111_0011_000: DATA = 1'b0;
            15'b10100111_0011_001: DATA = 1'b0;
            15'b10100111_0011_010: DATA = 1'b0;
            15'b10100111_0011_011: DATA = 1'b0;
            15'b10100111_0011_100: DATA = 1'b0;
            15'b10100111_0011_101: DATA = 1'b0;
            15'b10100111_0011_110: DATA = 1'b0;
            15'b10100111_0011_111: DATA = 1'b1;
            // SQUARE- ROW 1 COL 4 Row 4
            15'b10100111_0100_000: DATA = 1'b0;
            15'b10100111_0100_001: DATA = 1'b0;
            15'b10100111_0100_010: DATA = 1'b0;
            15'b10100111_0100_011: DATA = 1'b0;
            15'b10100111_0100_100: DATA = 1'b0;
            15'b10100111_0100_101: DATA = 1'b0;
            15'b10100111_0100_110: DATA = 1'b0;
            15'b10100111_0100_111: DATA = 1'b1;
            // SQUARE- ROW 1 COL 4 Row 5
            15'b10100111_0101_000: DATA = 1'b0;
            15'b10100111_0101_001: DATA = 1'b0;
            15'b10100111_0101_010: DATA = 1'b0;
            15'b10100111_0101_011: DATA = 1'b0;
            15'b10100111_0101_100: DATA = 1'b0;
            15'b10100111_0101_101: DATA = 1'b0;
            15'b10100111_0101_110: DATA = 1'b0;
            15'b10100111_0101_111: DATA = 1'b1;
            // SQUARE- ROW 1 COL 4 Row 6
            15'b10100111_0110_000: DATA = 1'b0;
            15'b10100111_0110_001: DATA = 1'b0;
            15'b10100111_0110_010: DATA = 1'b0;
            15'b10100111_0110_011: DATA = 1'b0;
            15'b10100111_0110_100: DATA = 1'b0;
            15'b10100111_0110_101: DATA = 1'b0;
            15'b10100111_0110_110: DATA = 1'b0;
            15'b10100111_0110_111: DATA = 1'b1;
            // SQUARE- ROW 1 COL 4 Row 7
            15'b10100111_0111_000: DATA = 1'b0;
            15'b10100111_0111_001: DATA = 1'b0;
            15'b10100111_0111_010: DATA = 1'b0;
            15'b10100111_0111_011: DATA = 1'b0;
            15'b10100111_0111_100: DATA = 1'b0;
            15'b10100111_0111_101: DATA = 1'b0;
            15'b10100111_0111_110: DATA = 1'b0;
            15'b10100111_0111_111: DATA = 1'b1;
            // SQUARE- ROW 1 COL 4 Row 8
            15'b10100111_1000_000: DATA = 1'b0;
            15'b10100111_1000_001: DATA = 1'b0;
            15'b10100111_1000_010: DATA = 1'b0;
            15'b10100111_1000_011: DATA = 1'b0;
            15'b10100111_1000_100: DATA = 1'b0;
            15'b10100111_1000_101: DATA = 1'b0;
            15'b10100111_1000_110: DATA = 1'b0;
            15'b10100111_1000_111: DATA = 1'b1;
            // SQUARE- ROW 1 COL 4 Row 9
            15'b10100111_1001_000: DATA = 1'b0;
            15'b10100111_1001_001: DATA = 1'b0;
            15'b10100111_1001_010: DATA = 1'b0;
            15'b10100111_1001_011: DATA = 1'b0;
            15'b10100111_1001_100: DATA = 1'b0;
            15'b10100111_1001_101: DATA = 1'b0;
            15'b10100111_1001_110: DATA = 1'b0;
            15'b10100111_1001_111: DATA = 1'b1;
            // SQUARE- ROW 1 COL 4 Row 10
            15'b10100111_1010_000: DATA = 1'b0;
            15'b10100111_1010_001: DATA = 1'b0;
            15'b10100111_1010_010: DATA = 1'b0;
            15'b10100111_1010_011: DATA = 1'b0;
            15'b10100111_1010_100: DATA = 1'b0;
            15'b10100111_1010_101: DATA = 1'b0;
            15'b10100111_1010_110: DATA = 1'b0;
            15'b10100111_1010_111: DATA = 1'b1;
            // SQUARE- ROW 1 COL 4 Row 11
            15'b10100111_1011_000: DATA = 1'b0;
            15'b10100111_1011_001: DATA = 1'b0;
            15'b10100111_1011_010: DATA = 1'b0;
            15'b10100111_1011_011: DATA = 1'b0;
            15'b10100111_1011_100: DATA = 1'b0;
            15'b10100111_1011_101: DATA = 1'b0;
            15'b10100111_1011_110: DATA = 1'b0;
            15'b10100111_1011_111: DATA = 1'b1;
            // SQUARE- ROW 1 COL 4 Row 12
            15'b10100111_1100_000: DATA = 1'b0;
            15'b10100111_1100_001: DATA = 1'b0;
            15'b10100111_1100_010: DATA = 1'b0;
            15'b10100111_1100_011: DATA = 1'b0;
            15'b10100111_1100_100: DATA = 1'b0;
            15'b10100111_1100_101: DATA = 1'b0;
            15'b10100111_1100_110: DATA = 1'b0;
            15'b10100111_1100_111: DATA = 1'b1;
            // SQUARE- ROW 1 COL 4 Row 13
            15'b10100111_1101_000: DATA = 1'b0;
            15'b10100111_1101_001: DATA = 1'b0;
            15'b10100111_1101_010: DATA = 1'b0;
            15'b10100111_1101_011: DATA = 1'b0;
            15'b10100111_1101_100: DATA = 1'b0;
            15'b10100111_1101_101: DATA = 1'b0;
            15'b10100111_1101_110: DATA = 1'b0;
            15'b10100111_1101_111: DATA = 1'b1;
            // SQUARE- ROW 1 COL 4 Row 14
            15'b10100111_1110_000: DATA = 1'b0;
            15'b10100111_1110_001: DATA = 1'b0;
            15'b10100111_1110_010: DATA = 1'b0;
            15'b10100111_1110_011: DATA = 1'b0;
            15'b10100111_1110_100: DATA = 1'b0;
            15'b10100111_1110_101: DATA = 1'b0;
            15'b10100111_1110_110: DATA = 1'b0;
            15'b10100111_1110_111: DATA = 1'b1;
            // SQUARE- ROW 1 COL 4 Row 15
            15'b10100111_1111_000: DATA = 1'b1;
            15'b10100111_1111_001: DATA = 1'b1;
            15'b10100111_1111_010: DATA = 1'b1;
            15'b10100111_1111_011: DATA = 1'b1;
            15'b10100111_1111_100: DATA = 1'b1;
            15'b10100111_1111_101: DATA = 1'b1;
            15'b10100111_1111_110: DATA = 1'b1;
            15'b10100111_1111_111: DATA = 1'b1;
            // TRIANGLE+ ROW 0 COL 0 Row 0
            15'b10101000_0000_000: DATA = 1'b0;
            15'b10101000_0000_001: DATA = 1'b0;
            15'b10101000_0000_010: DATA = 1'b0;
            15'b10101000_0000_011: DATA = 1'b0;
            15'b10101000_0000_100: DATA = 1'b0;
            15'b10101000_0000_101: DATA = 1'b0;
            15'b10101000_0000_110: DATA = 1'b0;
            15'b10101000_0000_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 0 Row 1
            15'b10101000_0001_000: DATA = 1'b0;
            15'b10101000_0001_001: DATA = 1'b0;
            15'b10101000_0001_010: DATA = 1'b0;
            15'b10101000_0001_011: DATA = 1'b0;
            15'b10101000_0001_100: DATA = 1'b0;
            15'b10101000_0001_101: DATA = 1'b0;
            15'b10101000_0001_110: DATA = 1'b0;
            15'b10101000_0001_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 0 Row 2
            15'b10101000_0010_000: DATA = 1'b0;
            15'b10101000_0010_001: DATA = 1'b0;
            15'b10101000_0010_010: DATA = 1'b0;
            15'b10101000_0010_011: DATA = 1'b0;
            15'b10101000_0010_100: DATA = 1'b0;
            15'b10101000_0010_101: DATA = 1'b0;
            15'b10101000_0010_110: DATA = 1'b0;
            15'b10101000_0010_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 0 Row 3
            15'b10101000_0011_000: DATA = 1'b0;
            15'b10101000_0011_001: DATA = 1'b0;
            15'b10101000_0011_010: DATA = 1'b0;
            15'b10101000_0011_011: DATA = 1'b0;
            15'b10101000_0011_100: DATA = 1'b0;
            15'b10101000_0011_101: DATA = 1'b0;
            15'b10101000_0011_110: DATA = 1'b0;
            15'b10101000_0011_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 0 Row 4
            15'b10101000_0100_000: DATA = 1'b0;
            15'b10101000_0100_001: DATA = 1'b0;
            15'b10101000_0100_010: DATA = 1'b0;
            15'b10101000_0100_011: DATA = 1'b0;
            15'b10101000_0100_100: DATA = 1'b0;
            15'b10101000_0100_101: DATA = 1'b0;
            15'b10101000_0100_110: DATA = 1'b0;
            15'b10101000_0100_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 0 Row 5
            15'b10101000_0101_000: DATA = 1'b0;
            15'b10101000_0101_001: DATA = 1'b0;
            15'b10101000_0101_010: DATA = 1'b0;
            15'b10101000_0101_011: DATA = 1'b0;
            15'b10101000_0101_100: DATA = 1'b0;
            15'b10101000_0101_101: DATA = 1'b0;
            15'b10101000_0101_110: DATA = 1'b0;
            15'b10101000_0101_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 0 Row 6
            15'b10101000_0110_000: DATA = 1'b0;
            15'b10101000_0110_001: DATA = 1'b0;
            15'b10101000_0110_010: DATA = 1'b0;
            15'b10101000_0110_011: DATA = 1'b0;
            15'b10101000_0110_100: DATA = 1'b0;
            15'b10101000_0110_101: DATA = 1'b0;
            15'b10101000_0110_110: DATA = 1'b0;
            15'b10101000_0110_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 0 Row 7
            15'b10101000_0111_000: DATA = 1'b0;
            15'b10101000_0111_001: DATA = 1'b0;
            15'b10101000_0111_010: DATA = 1'b0;
            15'b10101000_0111_011: DATA = 1'b0;
            15'b10101000_0111_100: DATA = 1'b0;
            15'b10101000_0111_101: DATA = 1'b0;
            15'b10101000_0111_110: DATA = 1'b0;
            15'b10101000_0111_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 0 Row 8
            15'b10101000_1000_000: DATA = 1'b0;
            15'b10101000_1000_001: DATA = 1'b0;
            15'b10101000_1000_010: DATA = 1'b0;
            15'b10101000_1000_011: DATA = 1'b0;
            15'b10101000_1000_100: DATA = 1'b0;
            15'b10101000_1000_101: DATA = 1'b0;
            15'b10101000_1000_110: DATA = 1'b0;
            15'b10101000_1000_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 0 Row 9
            15'b10101000_1001_000: DATA = 1'b0;
            15'b10101000_1001_001: DATA = 1'b0;
            15'b10101000_1001_010: DATA = 1'b0;
            15'b10101000_1001_011: DATA = 1'b0;
            15'b10101000_1001_100: DATA = 1'b0;
            15'b10101000_1001_101: DATA = 1'b0;
            15'b10101000_1001_110: DATA = 1'b0;
            15'b10101000_1001_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 0 Row 10
            15'b10101000_1010_000: DATA = 1'b0;
            15'b10101000_1010_001: DATA = 1'b0;
            15'b10101000_1010_010: DATA = 1'b0;
            15'b10101000_1010_011: DATA = 1'b0;
            15'b10101000_1010_100: DATA = 1'b0;
            15'b10101000_1010_101: DATA = 1'b0;
            15'b10101000_1010_110: DATA = 1'b0;
            15'b10101000_1010_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 0 Row 11
            15'b10101000_1011_000: DATA = 1'b0;
            15'b10101000_1011_001: DATA = 1'b0;
            15'b10101000_1011_010: DATA = 1'b0;
            15'b10101000_1011_011: DATA = 1'b0;
            15'b10101000_1011_100: DATA = 1'b0;
            15'b10101000_1011_101: DATA = 1'b0;
            15'b10101000_1011_110: DATA = 1'b0;
            15'b10101000_1011_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 0 Row 12
            15'b10101000_1100_000: DATA = 1'b0;
            15'b10101000_1100_001: DATA = 1'b0;
            15'b10101000_1100_010: DATA = 1'b0;
            15'b10101000_1100_011: DATA = 1'b0;
            15'b10101000_1100_100: DATA = 1'b0;
            15'b10101000_1100_101: DATA = 1'b0;
            15'b10101000_1100_110: DATA = 1'b0;
            15'b10101000_1100_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 0 Row 13
            15'b10101000_1101_000: DATA = 1'b0;
            15'b10101000_1101_001: DATA = 1'b0;
            15'b10101000_1101_010: DATA = 1'b0;
            15'b10101000_1101_011: DATA = 1'b0;
            15'b10101000_1101_100: DATA = 1'b0;
            15'b10101000_1101_101: DATA = 1'b0;
            15'b10101000_1101_110: DATA = 1'b0;
            15'b10101000_1101_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 0 Row 14
            15'b10101000_1110_000: DATA = 1'b0;
            15'b10101000_1110_001: DATA = 1'b0;
            15'b10101000_1110_010: DATA = 1'b0;
            15'b10101000_1110_011: DATA = 1'b0;
            15'b10101000_1110_100: DATA = 1'b0;
            15'b10101000_1110_101: DATA = 1'b0;
            15'b10101000_1110_110: DATA = 1'b0;
            15'b10101000_1110_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 0 Row 15
            15'b10101000_1111_000: DATA = 1'b0;
            15'b10101000_1111_001: DATA = 1'b0;
            15'b10101000_1111_010: DATA = 1'b0;
            15'b10101000_1111_011: DATA = 1'b0;
            15'b10101000_1111_100: DATA = 1'b0;
            15'b10101000_1111_101: DATA = 1'b0;
            15'b10101000_1111_110: DATA = 1'b0;
            15'b10101000_1111_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 1 Row 0
            15'b10101001_0000_000: DATA = 1'b0;
            15'b10101001_0000_001: DATA = 1'b0;
            15'b10101001_0000_010: DATA = 1'b0;
            15'b10101001_0000_011: DATA = 1'b0;
            15'b10101001_0000_100: DATA = 1'b0;
            15'b10101001_0000_101: DATA = 1'b0;
            15'b10101001_0000_110: DATA = 1'b0;
            15'b10101001_0000_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 1 Row 1
            15'b10101001_0001_000: DATA = 1'b0;
            15'b10101001_0001_001: DATA = 1'b0;
            15'b10101001_0001_010: DATA = 1'b0;
            15'b10101001_0001_011: DATA = 1'b0;
            15'b10101001_0001_100: DATA = 1'b0;
            15'b10101001_0001_101: DATA = 1'b0;
            15'b10101001_0001_110: DATA = 1'b0;
            15'b10101001_0001_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 1 Row 2
            15'b10101001_0010_000: DATA = 1'b0;
            15'b10101001_0010_001: DATA = 1'b0;
            15'b10101001_0010_010: DATA = 1'b0;
            15'b10101001_0010_011: DATA = 1'b0;
            15'b10101001_0010_100: DATA = 1'b0;
            15'b10101001_0010_101: DATA = 1'b0;
            15'b10101001_0010_110: DATA = 1'b0;
            15'b10101001_0010_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 1 Row 3
            15'b10101001_0011_000: DATA = 1'b0;
            15'b10101001_0011_001: DATA = 1'b0;
            15'b10101001_0011_010: DATA = 1'b0;
            15'b10101001_0011_011: DATA = 1'b0;
            15'b10101001_0011_100: DATA = 1'b0;
            15'b10101001_0011_101: DATA = 1'b0;
            15'b10101001_0011_110: DATA = 1'b0;
            15'b10101001_0011_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 1 Row 4
            15'b10101001_0100_000: DATA = 1'b0;
            15'b10101001_0100_001: DATA = 1'b0;
            15'b10101001_0100_010: DATA = 1'b0;
            15'b10101001_0100_011: DATA = 1'b0;
            15'b10101001_0100_100: DATA = 1'b0;
            15'b10101001_0100_101: DATA = 1'b0;
            15'b10101001_0100_110: DATA = 1'b0;
            15'b10101001_0100_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 1 Row 5
            15'b10101001_0101_000: DATA = 1'b0;
            15'b10101001_0101_001: DATA = 1'b0;
            15'b10101001_0101_010: DATA = 1'b0;
            15'b10101001_0101_011: DATA = 1'b0;
            15'b10101001_0101_100: DATA = 1'b0;
            15'b10101001_0101_101: DATA = 1'b0;
            15'b10101001_0101_110: DATA = 1'b0;
            15'b10101001_0101_111: DATA = 1'b1;
            // TRIANGLE+ ROW 0 COL 1 Row 6
            15'b10101001_0110_000: DATA = 1'b0;
            15'b10101001_0110_001: DATA = 1'b0;
            15'b10101001_0110_010: DATA = 1'b0;
            15'b10101001_0110_011: DATA = 1'b0;
            15'b10101001_0110_100: DATA = 1'b0;
            15'b10101001_0110_101: DATA = 1'b0;
            15'b10101001_0110_110: DATA = 1'b1;
            15'b10101001_0110_111: DATA = 1'b1;
            // TRIANGLE+ ROW 0 COL 1 Row 7
            15'b10101001_0111_000: DATA = 1'b0;
            15'b10101001_0111_001: DATA = 1'b0;
            15'b10101001_0111_010: DATA = 1'b0;
            15'b10101001_0111_011: DATA = 1'b0;
            15'b10101001_0111_100: DATA = 1'b0;
            15'b10101001_0111_101: DATA = 1'b0;
            15'b10101001_0111_110: DATA = 1'b1;
            15'b10101001_0111_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 1 Row 8
            15'b10101001_1000_000: DATA = 1'b0;
            15'b10101001_1000_001: DATA = 1'b0;
            15'b10101001_1000_010: DATA = 1'b0;
            15'b10101001_1000_011: DATA = 1'b0;
            15'b10101001_1000_100: DATA = 1'b0;
            15'b10101001_1000_101: DATA = 1'b1;
            15'b10101001_1000_110: DATA = 1'b1;
            15'b10101001_1000_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 1 Row 9
            15'b10101001_1001_000: DATA = 1'b0;
            15'b10101001_1001_001: DATA = 1'b0;
            15'b10101001_1001_010: DATA = 1'b0;
            15'b10101001_1001_011: DATA = 1'b0;
            15'b10101001_1001_100: DATA = 1'b0;
            15'b10101001_1001_101: DATA = 1'b1;
            15'b10101001_1001_110: DATA = 1'b0;
            15'b10101001_1001_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 1 Row 10
            15'b10101001_1010_000: DATA = 1'b0;
            15'b10101001_1010_001: DATA = 1'b0;
            15'b10101001_1010_010: DATA = 1'b0;
            15'b10101001_1010_011: DATA = 1'b0;
            15'b10101001_1010_100: DATA = 1'b1;
            15'b10101001_1010_101: DATA = 1'b1;
            15'b10101001_1010_110: DATA = 1'b0;
            15'b10101001_1010_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 1 Row 11
            15'b10101001_1011_000: DATA = 1'b0;
            15'b10101001_1011_001: DATA = 1'b0;
            15'b10101001_1011_010: DATA = 1'b0;
            15'b10101001_1011_011: DATA = 1'b1;
            15'b10101001_1011_100: DATA = 1'b1;
            15'b10101001_1011_101: DATA = 1'b0;
            15'b10101001_1011_110: DATA = 1'b0;
            15'b10101001_1011_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 1 Row 12
            15'b10101001_1100_000: DATA = 1'b0;
            15'b10101001_1100_001: DATA = 1'b0;
            15'b10101001_1100_010: DATA = 1'b0;
            15'b10101001_1100_011: DATA = 1'b1;
            15'b10101001_1100_100: DATA = 1'b0;
            15'b10101001_1100_101: DATA = 1'b0;
            15'b10101001_1100_110: DATA = 1'b0;
            15'b10101001_1100_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 1 Row 13
            15'b10101001_1101_000: DATA = 1'b0;
            15'b10101001_1101_001: DATA = 1'b0;
            15'b10101001_1101_010: DATA = 1'b1;
            15'b10101001_1101_011: DATA = 1'b1;
            15'b10101001_1101_100: DATA = 1'b0;
            15'b10101001_1101_101: DATA = 1'b0;
            15'b10101001_1101_110: DATA = 1'b0;
            15'b10101001_1101_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 1 Row 14
            15'b10101001_1110_000: DATA = 1'b0;
            15'b10101001_1110_001: DATA = 1'b0;
            15'b10101001_1110_010: DATA = 1'b1;
            15'b10101001_1110_011: DATA = 1'b0;
            15'b10101001_1110_100: DATA = 1'b0;
            15'b10101001_1110_101: DATA = 1'b0;
            15'b10101001_1110_110: DATA = 1'b0;
            15'b10101001_1110_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 1 Row 15
            15'b10101001_1111_000: DATA = 1'b0;
            15'b10101001_1111_001: DATA = 1'b1;
            15'b10101001_1111_010: DATA = 1'b1;
            15'b10101001_1111_011: DATA = 1'b0;
            15'b10101001_1111_100: DATA = 1'b0;
            15'b10101001_1111_101: DATA = 1'b0;
            15'b10101001_1111_110: DATA = 1'b0;
            15'b10101001_1111_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 2 Row 0
            15'b10101010_0000_000: DATA = 1'b0;
            15'b10101010_0000_001: DATA = 1'b0;
            15'b10101010_0000_010: DATA = 1'b0;
            15'b10101010_0000_011: DATA = 1'b1;
            15'b10101010_0000_100: DATA = 1'b1;
            15'b10101010_0000_101: DATA = 1'b0;
            15'b10101010_0000_110: DATA = 1'b0;
            15'b10101010_0000_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 2 Row 1
            15'b10101010_0001_000: DATA = 1'b0;
            15'b10101010_0001_001: DATA = 1'b1;
            15'b10101010_0001_010: DATA = 1'b1;
            15'b10101010_0001_011: DATA = 1'b0;
            15'b10101010_0001_100: DATA = 1'b0;
            15'b10101010_0001_101: DATA = 1'b1;
            15'b10101010_0001_110: DATA = 1'b1;
            15'b10101010_0001_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 2 Row 2
            15'b10101010_0010_000: DATA = 1'b0;
            15'b10101010_0010_001: DATA = 1'b1;
            15'b10101010_0010_010: DATA = 1'b0;
            15'b10101010_0010_011: DATA = 1'b0;
            15'b10101010_0010_100: DATA = 1'b0;
            15'b10101010_0010_101: DATA = 1'b0;
            15'b10101010_0010_110: DATA = 1'b1;
            15'b10101010_0010_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 2 Row 3
            15'b10101010_0011_000: DATA = 1'b1;
            15'b10101010_0011_001: DATA = 1'b1;
            15'b10101010_0011_010: DATA = 1'b0;
            15'b10101010_0011_011: DATA = 1'b0;
            15'b10101010_0011_100: DATA = 1'b0;
            15'b10101010_0011_101: DATA = 1'b0;
            15'b10101010_0011_110: DATA = 1'b1;
            15'b10101010_0011_111: DATA = 1'b1;
            // TRIANGLE+ ROW 0 COL 2 Row 4
            15'b10101010_0100_000: DATA = 1'b1;
            15'b10101010_0100_001: DATA = 1'b0;
            15'b10101010_0100_010: DATA = 1'b0;
            15'b10101010_0100_011: DATA = 1'b0;
            15'b10101010_0100_100: DATA = 1'b0;
            15'b10101010_0100_101: DATA = 1'b0;
            15'b10101010_0100_110: DATA = 1'b0;
            15'b10101010_0100_111: DATA = 1'b1;
            // TRIANGLE+ ROW 0 COL 2 Row 5
            15'b10101010_0101_000: DATA = 1'b1;
            15'b10101010_0101_001: DATA = 1'b0;
            15'b10101010_0101_010: DATA = 1'b0;
            15'b10101010_0101_011: DATA = 1'b0;
            15'b10101010_0101_100: DATA = 1'b0;
            15'b10101010_0101_101: DATA = 1'b0;
            15'b10101010_0101_110: DATA = 1'b0;
            15'b10101010_0101_111: DATA = 1'b1;
            // TRIANGLE+ ROW 0 COL 2 Row 6
            15'b10101010_0110_000: DATA = 1'b0;
            15'b10101010_0110_001: DATA = 1'b0;
            15'b10101010_0110_010: DATA = 1'b0;
            15'b10101010_0110_011: DATA = 1'b0;
            15'b10101010_0110_100: DATA = 1'b0;
            15'b10101010_0110_101: DATA = 1'b0;
            15'b10101010_0110_110: DATA = 1'b0;
            15'b10101010_0110_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 2 Row 7
            15'b10101010_0111_000: DATA = 1'b0;
            15'b10101010_0111_001: DATA = 1'b0;
            15'b10101010_0111_010: DATA = 1'b0;
            15'b10101010_0111_011: DATA = 1'b0;
            15'b10101010_0111_100: DATA = 1'b0;
            15'b10101010_0111_101: DATA = 1'b0;
            15'b10101010_0111_110: DATA = 1'b0;
            15'b10101010_0111_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 2 Row 8
            15'b10101010_1000_000: DATA = 1'b0;
            15'b10101010_1000_001: DATA = 1'b0;
            15'b10101010_1000_010: DATA = 1'b0;
            15'b10101010_1000_011: DATA = 1'b0;
            15'b10101010_1000_100: DATA = 1'b0;
            15'b10101010_1000_101: DATA = 1'b0;
            15'b10101010_1000_110: DATA = 1'b0;
            15'b10101010_1000_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 2 Row 9
            15'b10101010_1001_000: DATA = 1'b0;
            15'b10101010_1001_001: DATA = 1'b0;
            15'b10101010_1001_010: DATA = 1'b0;
            15'b10101010_1001_011: DATA = 1'b0;
            15'b10101010_1001_100: DATA = 1'b0;
            15'b10101010_1001_101: DATA = 1'b0;
            15'b10101010_1001_110: DATA = 1'b0;
            15'b10101010_1001_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 2 Row 10
            15'b10101010_1010_000: DATA = 1'b0;
            15'b10101010_1010_001: DATA = 1'b0;
            15'b10101010_1010_010: DATA = 1'b0;
            15'b10101010_1010_011: DATA = 1'b0;
            15'b10101010_1010_100: DATA = 1'b0;
            15'b10101010_1010_101: DATA = 1'b0;
            15'b10101010_1010_110: DATA = 1'b0;
            15'b10101010_1010_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 2 Row 11
            15'b10101010_1011_000: DATA = 1'b0;
            15'b10101010_1011_001: DATA = 1'b0;
            15'b10101010_1011_010: DATA = 1'b0;
            15'b10101010_1011_011: DATA = 1'b0;
            15'b10101010_1011_100: DATA = 1'b0;
            15'b10101010_1011_101: DATA = 1'b0;
            15'b10101010_1011_110: DATA = 1'b0;
            15'b10101010_1011_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 2 Row 12
            15'b10101010_1100_000: DATA = 1'b0;
            15'b10101010_1100_001: DATA = 1'b0;
            15'b10101010_1100_010: DATA = 1'b0;
            15'b10101010_1100_011: DATA = 1'b0;
            15'b10101010_1100_100: DATA = 1'b0;
            15'b10101010_1100_101: DATA = 1'b0;
            15'b10101010_1100_110: DATA = 1'b0;
            15'b10101010_1100_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 2 Row 13
            15'b10101010_1101_000: DATA = 1'b0;
            15'b10101010_1101_001: DATA = 1'b0;
            15'b10101010_1101_010: DATA = 1'b0;
            15'b10101010_1101_011: DATA = 1'b0;
            15'b10101010_1101_100: DATA = 1'b0;
            15'b10101010_1101_101: DATA = 1'b0;
            15'b10101010_1101_110: DATA = 1'b0;
            15'b10101010_1101_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 2 Row 14
            15'b10101010_1110_000: DATA = 1'b0;
            15'b10101010_1110_001: DATA = 1'b0;
            15'b10101010_1110_010: DATA = 1'b0;
            15'b10101010_1110_011: DATA = 1'b0;
            15'b10101010_1110_100: DATA = 1'b0;
            15'b10101010_1110_101: DATA = 1'b0;
            15'b10101010_1110_110: DATA = 1'b0;
            15'b10101010_1110_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 2 Row 15
            15'b10101010_1111_000: DATA = 1'b0;
            15'b10101010_1111_001: DATA = 1'b0;
            15'b10101010_1111_010: DATA = 1'b0;
            15'b10101010_1111_011: DATA = 1'b0;
            15'b10101010_1111_100: DATA = 1'b0;
            15'b10101010_1111_101: DATA = 1'b0;
            15'b10101010_1111_110: DATA = 1'b0;
            15'b10101010_1111_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 3 Row 0
            15'b10101011_0000_000: DATA = 1'b0;
            15'b10101011_0000_001: DATA = 1'b0;
            15'b10101011_0000_010: DATA = 1'b0;
            15'b10101011_0000_011: DATA = 1'b0;
            15'b10101011_0000_100: DATA = 1'b0;
            15'b10101011_0000_101: DATA = 1'b0;
            15'b10101011_0000_110: DATA = 1'b0;
            15'b10101011_0000_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 3 Row 1
            15'b10101011_0001_000: DATA = 1'b0;
            15'b10101011_0001_001: DATA = 1'b0;
            15'b10101011_0001_010: DATA = 1'b0;
            15'b10101011_0001_011: DATA = 1'b0;
            15'b10101011_0001_100: DATA = 1'b0;
            15'b10101011_0001_101: DATA = 1'b0;
            15'b10101011_0001_110: DATA = 1'b0;
            15'b10101011_0001_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 3 Row 2
            15'b10101011_0010_000: DATA = 1'b0;
            15'b10101011_0010_001: DATA = 1'b0;
            15'b10101011_0010_010: DATA = 1'b0;
            15'b10101011_0010_011: DATA = 1'b0;
            15'b10101011_0010_100: DATA = 1'b0;
            15'b10101011_0010_101: DATA = 1'b0;
            15'b10101011_0010_110: DATA = 1'b0;
            15'b10101011_0010_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 3 Row 3
            15'b10101011_0011_000: DATA = 1'b0;
            15'b10101011_0011_001: DATA = 1'b0;
            15'b10101011_0011_010: DATA = 1'b0;
            15'b10101011_0011_011: DATA = 1'b0;
            15'b10101011_0011_100: DATA = 1'b0;
            15'b10101011_0011_101: DATA = 1'b0;
            15'b10101011_0011_110: DATA = 1'b0;
            15'b10101011_0011_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 3 Row 4
            15'b10101011_0100_000: DATA = 1'b0;
            15'b10101011_0100_001: DATA = 1'b0;
            15'b10101011_0100_010: DATA = 1'b0;
            15'b10101011_0100_011: DATA = 1'b0;
            15'b10101011_0100_100: DATA = 1'b0;
            15'b10101011_0100_101: DATA = 1'b0;
            15'b10101011_0100_110: DATA = 1'b0;
            15'b10101011_0100_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 3 Row 5
            15'b10101011_0101_000: DATA = 1'b1;
            15'b10101011_0101_001: DATA = 1'b0;
            15'b10101011_0101_010: DATA = 1'b0;
            15'b10101011_0101_011: DATA = 1'b0;
            15'b10101011_0101_100: DATA = 1'b0;
            15'b10101011_0101_101: DATA = 1'b0;
            15'b10101011_0101_110: DATA = 1'b0;
            15'b10101011_0101_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 3 Row 6
            15'b10101011_0110_000: DATA = 1'b1;
            15'b10101011_0110_001: DATA = 1'b1;
            15'b10101011_0110_010: DATA = 1'b0;
            15'b10101011_0110_011: DATA = 1'b0;
            15'b10101011_0110_100: DATA = 1'b0;
            15'b10101011_0110_101: DATA = 1'b0;
            15'b10101011_0110_110: DATA = 1'b0;
            15'b10101011_0110_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 3 Row 7
            15'b10101011_0111_000: DATA = 1'b0;
            15'b10101011_0111_001: DATA = 1'b1;
            15'b10101011_0111_010: DATA = 1'b0;
            15'b10101011_0111_011: DATA = 1'b0;
            15'b10101011_0111_100: DATA = 1'b0;
            15'b10101011_0111_101: DATA = 1'b0;
            15'b10101011_0111_110: DATA = 1'b0;
            15'b10101011_0111_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 3 Row 8
            15'b10101011_1000_000: DATA = 1'b0;
            15'b10101011_1000_001: DATA = 1'b1;
            15'b10101011_1000_010: DATA = 1'b1;
            15'b10101011_1000_011: DATA = 1'b0;
            15'b10101011_1000_100: DATA = 1'b0;
            15'b10101011_1000_101: DATA = 1'b0;
            15'b10101011_1000_110: DATA = 1'b0;
            15'b10101011_1000_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 3 Row 9
            15'b10101011_1001_000: DATA = 1'b0;
            15'b10101011_1001_001: DATA = 1'b0;
            15'b10101011_1001_010: DATA = 1'b1;
            15'b10101011_1001_011: DATA = 1'b0;
            15'b10101011_1001_100: DATA = 1'b0;
            15'b10101011_1001_101: DATA = 1'b0;
            15'b10101011_1001_110: DATA = 1'b0;
            15'b10101011_1001_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 3 Row 10
            15'b10101011_1010_000: DATA = 1'b0;
            15'b10101011_1010_001: DATA = 1'b0;
            15'b10101011_1010_010: DATA = 1'b1;
            15'b10101011_1010_011: DATA = 1'b1;
            15'b10101011_1010_100: DATA = 1'b0;
            15'b10101011_1010_101: DATA = 1'b0;
            15'b10101011_1010_110: DATA = 1'b0;
            15'b10101011_1010_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 3 Row 11
            15'b10101011_1011_000: DATA = 1'b0;
            15'b10101011_1011_001: DATA = 1'b0;
            15'b10101011_1011_010: DATA = 1'b0;
            15'b10101011_1011_011: DATA = 1'b1;
            15'b10101011_1011_100: DATA = 1'b1;
            15'b10101011_1011_101: DATA = 1'b0;
            15'b10101011_1011_110: DATA = 1'b0;
            15'b10101011_1011_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 3 Row 12
            15'b10101011_1100_000: DATA = 1'b0;
            15'b10101011_1100_001: DATA = 1'b0;
            15'b10101011_1100_010: DATA = 1'b0;
            15'b10101011_1100_011: DATA = 1'b0;
            15'b10101011_1100_100: DATA = 1'b1;
            15'b10101011_1100_101: DATA = 1'b0;
            15'b10101011_1100_110: DATA = 1'b0;
            15'b10101011_1100_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 3 Row 13
            15'b10101011_1101_000: DATA = 1'b0;
            15'b10101011_1101_001: DATA = 1'b0;
            15'b10101011_1101_010: DATA = 1'b0;
            15'b10101011_1101_011: DATA = 1'b0;
            15'b10101011_1101_100: DATA = 1'b1;
            15'b10101011_1101_101: DATA = 1'b1;
            15'b10101011_1101_110: DATA = 1'b0;
            15'b10101011_1101_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 3 Row 14
            15'b10101011_1110_000: DATA = 1'b0;
            15'b10101011_1110_001: DATA = 1'b0;
            15'b10101011_1110_010: DATA = 1'b0;
            15'b10101011_1110_011: DATA = 1'b0;
            15'b10101011_1110_100: DATA = 1'b0;
            15'b10101011_1110_101: DATA = 1'b1;
            15'b10101011_1110_110: DATA = 1'b0;
            15'b10101011_1110_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 3 Row 15
            15'b10101011_1111_000: DATA = 1'b0;
            15'b10101011_1111_001: DATA = 1'b0;
            15'b10101011_1111_010: DATA = 1'b0;
            15'b10101011_1111_011: DATA = 1'b0;
            15'b10101011_1111_100: DATA = 1'b0;
            15'b10101011_1111_101: DATA = 1'b1;
            15'b10101011_1111_110: DATA = 1'b1;
            15'b10101011_1111_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 4 Row 0
            15'b10101100_0000_000: DATA = 1'b0;
            15'b10101100_0000_001: DATA = 1'b0;
            15'b10101100_0000_010: DATA = 1'b0;
            15'b10101100_0000_011: DATA = 1'b0;
            15'b10101100_0000_100: DATA = 1'b0;
            15'b10101100_0000_101: DATA = 1'b0;
            15'b10101100_0000_110: DATA = 1'b0;
            15'b10101100_0000_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 4 Row 1
            15'b10101100_0001_000: DATA = 1'b0;
            15'b10101100_0001_001: DATA = 1'b0;
            15'b10101100_0001_010: DATA = 1'b0;
            15'b10101100_0001_011: DATA = 1'b0;
            15'b10101100_0001_100: DATA = 1'b0;
            15'b10101100_0001_101: DATA = 1'b0;
            15'b10101100_0001_110: DATA = 1'b0;
            15'b10101100_0001_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 4 Row 2
            15'b10101100_0010_000: DATA = 1'b0;
            15'b10101100_0010_001: DATA = 1'b0;
            15'b10101100_0010_010: DATA = 1'b0;
            15'b10101100_0010_011: DATA = 1'b0;
            15'b10101100_0010_100: DATA = 1'b0;
            15'b10101100_0010_101: DATA = 1'b0;
            15'b10101100_0010_110: DATA = 1'b0;
            15'b10101100_0010_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 4 Row 3
            15'b10101100_0011_000: DATA = 1'b0;
            15'b10101100_0011_001: DATA = 1'b0;
            15'b10101100_0011_010: DATA = 1'b0;
            15'b10101100_0011_011: DATA = 1'b0;
            15'b10101100_0011_100: DATA = 1'b0;
            15'b10101100_0011_101: DATA = 1'b0;
            15'b10101100_0011_110: DATA = 1'b0;
            15'b10101100_0011_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 4 Row 4
            15'b10101100_0100_000: DATA = 1'b0;
            15'b10101100_0100_001: DATA = 1'b0;
            15'b10101100_0100_010: DATA = 1'b0;
            15'b10101100_0100_011: DATA = 1'b0;
            15'b10101100_0100_100: DATA = 1'b0;
            15'b10101100_0100_101: DATA = 1'b0;
            15'b10101100_0100_110: DATA = 1'b0;
            15'b10101100_0100_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 4 Row 5
            15'b10101100_0101_000: DATA = 1'b0;
            15'b10101100_0101_001: DATA = 1'b0;
            15'b10101100_0101_010: DATA = 1'b0;
            15'b10101100_0101_011: DATA = 1'b0;
            15'b10101100_0101_100: DATA = 1'b0;
            15'b10101100_0101_101: DATA = 1'b0;
            15'b10101100_0101_110: DATA = 1'b0;
            15'b10101100_0101_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 4 Row 6
            15'b10101100_0110_000: DATA = 1'b0;
            15'b10101100_0110_001: DATA = 1'b0;
            15'b10101100_0110_010: DATA = 1'b0;
            15'b10101100_0110_011: DATA = 1'b0;
            15'b10101100_0110_100: DATA = 1'b0;
            15'b10101100_0110_101: DATA = 1'b0;
            15'b10101100_0110_110: DATA = 1'b0;
            15'b10101100_0110_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 4 Row 7
            15'b10101100_0111_000: DATA = 1'b0;
            15'b10101100_0111_001: DATA = 1'b0;
            15'b10101100_0111_010: DATA = 1'b0;
            15'b10101100_0111_011: DATA = 1'b0;
            15'b10101100_0111_100: DATA = 1'b0;
            15'b10101100_0111_101: DATA = 1'b0;
            15'b10101100_0111_110: DATA = 1'b0;
            15'b10101100_0111_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 4 Row 8
            15'b10101100_1000_000: DATA = 1'b0;
            15'b10101100_1000_001: DATA = 1'b0;
            15'b10101100_1000_010: DATA = 1'b0;
            15'b10101100_1000_011: DATA = 1'b0;
            15'b10101100_1000_100: DATA = 1'b0;
            15'b10101100_1000_101: DATA = 1'b0;
            15'b10101100_1000_110: DATA = 1'b0;
            15'b10101100_1000_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 4 Row 9
            15'b10101100_1001_000: DATA = 1'b0;
            15'b10101100_1001_001: DATA = 1'b0;
            15'b10101100_1001_010: DATA = 1'b0;
            15'b10101100_1001_011: DATA = 1'b0;
            15'b10101100_1001_100: DATA = 1'b0;
            15'b10101100_1001_101: DATA = 1'b0;
            15'b10101100_1001_110: DATA = 1'b0;
            15'b10101100_1001_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 4 Row 10
            15'b10101100_1010_000: DATA = 1'b0;
            15'b10101100_1010_001: DATA = 1'b0;
            15'b10101100_1010_010: DATA = 1'b0;
            15'b10101100_1010_011: DATA = 1'b0;
            15'b10101100_1010_100: DATA = 1'b0;
            15'b10101100_1010_101: DATA = 1'b0;
            15'b10101100_1010_110: DATA = 1'b0;
            15'b10101100_1010_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 4 Row 11
            15'b10101100_1011_000: DATA = 1'b0;
            15'b10101100_1011_001: DATA = 1'b0;
            15'b10101100_1011_010: DATA = 1'b0;
            15'b10101100_1011_011: DATA = 1'b0;
            15'b10101100_1011_100: DATA = 1'b0;
            15'b10101100_1011_101: DATA = 1'b0;
            15'b10101100_1011_110: DATA = 1'b0;
            15'b10101100_1011_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 4 Row 12
            15'b10101100_1100_000: DATA = 1'b0;
            15'b10101100_1100_001: DATA = 1'b0;
            15'b10101100_1100_010: DATA = 1'b0;
            15'b10101100_1100_011: DATA = 1'b0;
            15'b10101100_1100_100: DATA = 1'b0;
            15'b10101100_1100_101: DATA = 1'b0;
            15'b10101100_1100_110: DATA = 1'b0;
            15'b10101100_1100_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 4 Row 13
            15'b10101100_1101_000: DATA = 1'b0;
            15'b10101100_1101_001: DATA = 1'b0;
            15'b10101100_1101_010: DATA = 1'b0;
            15'b10101100_1101_011: DATA = 1'b0;
            15'b10101100_1101_100: DATA = 1'b0;
            15'b10101100_1101_101: DATA = 1'b0;
            15'b10101100_1101_110: DATA = 1'b0;
            15'b10101100_1101_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 4 Row 14
            15'b10101100_1110_000: DATA = 1'b0;
            15'b10101100_1110_001: DATA = 1'b0;
            15'b10101100_1110_010: DATA = 1'b0;
            15'b10101100_1110_011: DATA = 1'b0;
            15'b10101100_1110_100: DATA = 1'b0;
            15'b10101100_1110_101: DATA = 1'b0;
            15'b10101100_1110_110: DATA = 1'b0;
            15'b10101100_1110_111: DATA = 1'b0;
            // TRIANGLE+ ROW 0 COL 4 Row 15
            15'b10101100_1111_000: DATA = 1'b0;
            15'b10101100_1111_001: DATA = 1'b0;
            15'b10101100_1111_010: DATA = 1'b0;
            15'b10101100_1111_011: DATA = 1'b0;
            15'b10101100_1111_100: DATA = 1'b0;
            15'b10101100_1111_101: DATA = 1'b0;
            15'b10101100_1111_110: DATA = 1'b0;
            15'b10101100_1111_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 0 Row 0
            15'b10101101_0000_000: DATA = 1'b0;
            15'b10101101_0000_001: DATA = 1'b0;
            15'b10101101_0000_010: DATA = 1'b0;
            15'b10101101_0000_011: DATA = 1'b0;
            15'b10101101_0000_100: DATA = 1'b0;
            15'b10101101_0000_101: DATA = 1'b0;
            15'b10101101_0000_110: DATA = 1'b0;
            15'b10101101_0000_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 0 Row 1
            15'b10101101_0001_000: DATA = 1'b0;
            15'b10101101_0001_001: DATA = 1'b0;
            15'b10101101_0001_010: DATA = 1'b0;
            15'b10101101_0001_011: DATA = 1'b0;
            15'b10101101_0001_100: DATA = 1'b0;
            15'b10101101_0001_101: DATA = 1'b0;
            15'b10101101_0001_110: DATA = 1'b0;
            15'b10101101_0001_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 0 Row 2
            15'b10101101_0010_000: DATA = 1'b0;
            15'b10101101_0010_001: DATA = 1'b0;
            15'b10101101_0010_010: DATA = 1'b0;
            15'b10101101_0010_011: DATA = 1'b0;
            15'b10101101_0010_100: DATA = 1'b0;
            15'b10101101_0010_101: DATA = 1'b0;
            15'b10101101_0010_110: DATA = 1'b0;
            15'b10101101_0010_111: DATA = 1'b1;
            // TRIANGLE+ ROW 1 COL 0 Row 3
            15'b10101101_0011_000: DATA = 1'b0;
            15'b10101101_0011_001: DATA = 1'b0;
            15'b10101101_0011_010: DATA = 1'b0;
            15'b10101101_0011_011: DATA = 1'b0;
            15'b10101101_0011_100: DATA = 1'b0;
            15'b10101101_0011_101: DATA = 1'b0;
            15'b10101101_0011_110: DATA = 1'b0;
            15'b10101101_0011_111: DATA = 1'b1;
            // TRIANGLE+ ROW 1 COL 0 Row 4
            15'b10101101_0100_000: DATA = 1'b0;
            15'b10101101_0100_001: DATA = 1'b0;
            15'b10101101_0100_010: DATA = 1'b0;
            15'b10101101_0100_011: DATA = 1'b0;
            15'b10101101_0100_100: DATA = 1'b0;
            15'b10101101_0100_101: DATA = 1'b0;
            15'b10101101_0100_110: DATA = 1'b1;
            15'b10101101_0100_111: DATA = 1'b1;
            // TRIANGLE+ ROW 1 COL 0 Row 5
            15'b10101101_0101_000: DATA = 1'b0;
            15'b10101101_0101_001: DATA = 1'b0;
            15'b10101101_0101_010: DATA = 1'b0;
            15'b10101101_0101_011: DATA = 1'b0;
            15'b10101101_0101_100: DATA = 1'b0;
            15'b10101101_0101_101: DATA = 1'b1;
            15'b10101101_0101_110: DATA = 1'b1;
            15'b10101101_0101_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 0 Row 6
            15'b10101101_0110_000: DATA = 1'b0;
            15'b10101101_0110_001: DATA = 1'b0;
            15'b10101101_0110_010: DATA = 1'b0;
            15'b10101101_0110_011: DATA = 1'b0;
            15'b10101101_0110_100: DATA = 1'b0;
            15'b10101101_0110_101: DATA = 1'b1;
            15'b10101101_0110_110: DATA = 1'b0;
            15'b10101101_0110_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 0 Row 7
            15'b10101101_0111_000: DATA = 1'b0;
            15'b10101101_0111_001: DATA = 1'b0;
            15'b10101101_0111_010: DATA = 1'b0;
            15'b10101101_0111_011: DATA = 1'b0;
            15'b10101101_0111_100: DATA = 1'b1;
            15'b10101101_0111_101: DATA = 1'b1;
            15'b10101101_0111_110: DATA = 1'b0;
            15'b10101101_0111_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 0 Row 8
            15'b10101101_1000_000: DATA = 1'b0;
            15'b10101101_1000_001: DATA = 1'b0;
            15'b10101101_1000_010: DATA = 1'b0;
            15'b10101101_1000_011: DATA = 1'b0;
            15'b10101101_1000_100: DATA = 1'b1;
            15'b10101101_1000_101: DATA = 1'b0;
            15'b10101101_1000_110: DATA = 1'b0;
            15'b10101101_1000_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 0 Row 9
            15'b10101101_1001_000: DATA = 1'b0;
            15'b10101101_1001_001: DATA = 1'b0;
            15'b10101101_1001_010: DATA = 1'b0;
            15'b10101101_1001_011: DATA = 1'b1;
            15'b10101101_1001_100: DATA = 1'b1;
            15'b10101101_1001_101: DATA = 1'b0;
            15'b10101101_1001_110: DATA = 1'b0;
            15'b10101101_1001_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 0 Row 10
            15'b10101101_1010_000: DATA = 1'b0;
            15'b10101101_1010_001: DATA = 1'b0;
            15'b10101101_1010_010: DATA = 1'b1;
            15'b10101101_1010_011: DATA = 1'b1;
            15'b10101101_1010_100: DATA = 1'b0;
            15'b10101101_1010_101: DATA = 1'b0;
            15'b10101101_1010_110: DATA = 1'b0;
            15'b10101101_1010_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 0 Row 11
            15'b10101101_1011_000: DATA = 1'b0;
            15'b10101101_1011_001: DATA = 1'b0;
            15'b10101101_1011_010: DATA = 1'b1;
            15'b10101101_1011_011: DATA = 1'b0;
            15'b10101101_1011_100: DATA = 1'b0;
            15'b10101101_1011_101: DATA = 1'b0;
            15'b10101101_1011_110: DATA = 1'b0;
            15'b10101101_1011_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 0 Row 12
            15'b10101101_1100_000: DATA = 1'b0;
            15'b10101101_1100_001: DATA = 1'b1;
            15'b10101101_1100_010: DATA = 1'b1;
            15'b10101101_1100_011: DATA = 1'b0;
            15'b10101101_1100_100: DATA = 1'b0;
            15'b10101101_1100_101: DATA = 1'b0;
            15'b10101101_1100_110: DATA = 1'b0;
            15'b10101101_1100_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 0 Row 13
            15'b10101101_1101_000: DATA = 1'b0;
            15'b10101101_1101_001: DATA = 1'b1;
            15'b10101101_1101_010: DATA = 1'b0;
            15'b10101101_1101_011: DATA = 1'b0;
            15'b10101101_1101_100: DATA = 1'b0;
            15'b10101101_1101_101: DATA = 1'b0;
            15'b10101101_1101_110: DATA = 1'b0;
            15'b10101101_1101_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 0 Row 14
            15'b10101101_1110_000: DATA = 1'b1;
            15'b10101101_1110_001: DATA = 1'b1;
            15'b10101101_1110_010: DATA = 1'b0;
            15'b10101101_1110_011: DATA = 1'b0;
            15'b10101101_1110_100: DATA = 1'b0;
            15'b10101101_1110_101: DATA = 1'b0;
            15'b10101101_1110_110: DATA = 1'b0;
            15'b10101101_1110_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 0 Row 15
            15'b10101101_1111_000: DATA = 1'b1;
            15'b10101101_1111_001: DATA = 1'b0;
            15'b10101101_1111_010: DATA = 1'b0;
            15'b10101101_1111_011: DATA = 1'b0;
            15'b10101101_1111_100: DATA = 1'b0;
            15'b10101101_1111_101: DATA = 1'b0;
            15'b10101101_1111_110: DATA = 1'b0;
            15'b10101101_1111_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 1 Row 0
            15'b10101110_0000_000: DATA = 1'b1;
            15'b10101110_0000_001: DATA = 1'b1;
            15'b10101110_0000_010: DATA = 1'b0;
            15'b10101110_0000_011: DATA = 1'b0;
            15'b10101110_0000_100: DATA = 1'b0;
            15'b10101110_0000_101: DATA = 1'b0;
            15'b10101110_0000_110: DATA = 1'b0;
            15'b10101110_0000_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 1 Row 1
            15'b10101110_0001_000: DATA = 1'b1;
            15'b10101110_0001_001: DATA = 1'b0;
            15'b10101110_0001_010: DATA = 1'b0;
            15'b10101110_0001_011: DATA = 1'b0;
            15'b10101110_0001_100: DATA = 1'b0;
            15'b10101110_0001_101: DATA = 1'b0;
            15'b10101110_0001_110: DATA = 1'b0;
            15'b10101110_0001_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 1 Row 2
            15'b10101110_0010_000: DATA = 1'b1;
            15'b10101110_0010_001: DATA = 1'b0;
            15'b10101110_0010_010: DATA = 1'b0;
            15'b10101110_0010_011: DATA = 1'b0;
            15'b10101110_0010_100: DATA = 1'b0;
            15'b10101110_0010_101: DATA = 1'b0;
            15'b10101110_0010_110: DATA = 1'b0;
            15'b10101110_0010_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 1 Row 3
            15'b10101110_0011_000: DATA = 1'b0;
            15'b10101110_0011_001: DATA = 1'b0;
            15'b10101110_0011_010: DATA = 1'b0;
            15'b10101110_0011_011: DATA = 1'b0;
            15'b10101110_0011_100: DATA = 1'b0;
            15'b10101110_0011_101: DATA = 1'b0;
            15'b10101110_0011_110: DATA = 1'b0;
            15'b10101110_0011_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 1 Row 4
            15'b10101110_0100_000: DATA = 1'b0;
            15'b10101110_0100_001: DATA = 1'b0;
            15'b10101110_0100_010: DATA = 1'b0;
            15'b10101110_0100_011: DATA = 1'b0;
            15'b10101110_0100_100: DATA = 1'b0;
            15'b10101110_0100_101: DATA = 1'b0;
            15'b10101110_0100_110: DATA = 1'b0;
            15'b10101110_0100_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 1 Row 5
            15'b10101110_0101_000: DATA = 1'b0;
            15'b10101110_0101_001: DATA = 1'b0;
            15'b10101110_0101_010: DATA = 1'b0;
            15'b10101110_0101_011: DATA = 1'b0;
            15'b10101110_0101_100: DATA = 1'b0;
            15'b10101110_0101_101: DATA = 1'b0;
            15'b10101110_0101_110: DATA = 1'b0;
            15'b10101110_0101_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 1 Row 6
            15'b10101110_0110_000: DATA = 1'b0;
            15'b10101110_0110_001: DATA = 1'b0;
            15'b10101110_0110_010: DATA = 1'b0;
            15'b10101110_0110_011: DATA = 1'b0;
            15'b10101110_0110_100: DATA = 1'b0;
            15'b10101110_0110_101: DATA = 1'b0;
            15'b10101110_0110_110: DATA = 1'b0;
            15'b10101110_0110_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 1 Row 7
            15'b10101110_0111_000: DATA = 1'b0;
            15'b10101110_0111_001: DATA = 1'b0;
            15'b10101110_0111_010: DATA = 1'b0;
            15'b10101110_0111_011: DATA = 1'b0;
            15'b10101110_0111_100: DATA = 1'b0;
            15'b10101110_0111_101: DATA = 1'b0;
            15'b10101110_0111_110: DATA = 1'b0;
            15'b10101110_0111_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 1 Row 8
            15'b10101110_1000_000: DATA = 1'b0;
            15'b10101110_1000_001: DATA = 1'b0;
            15'b10101110_1000_010: DATA = 1'b0;
            15'b10101110_1000_011: DATA = 1'b0;
            15'b10101110_1000_100: DATA = 1'b0;
            15'b10101110_1000_101: DATA = 1'b0;
            15'b10101110_1000_110: DATA = 1'b0;
            15'b10101110_1000_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 1 Row 9
            15'b10101110_1001_000: DATA = 1'b0;
            15'b10101110_1001_001: DATA = 1'b0;
            15'b10101110_1001_010: DATA = 1'b0;
            15'b10101110_1001_011: DATA = 1'b0;
            15'b10101110_1001_100: DATA = 1'b0;
            15'b10101110_1001_101: DATA = 1'b0;
            15'b10101110_1001_110: DATA = 1'b0;
            15'b10101110_1001_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 1 Row 10
            15'b10101110_1010_000: DATA = 1'b0;
            15'b10101110_1010_001: DATA = 1'b0;
            15'b10101110_1010_010: DATA = 1'b0;
            15'b10101110_1010_011: DATA = 1'b0;
            15'b10101110_1010_100: DATA = 1'b0;
            15'b10101110_1010_101: DATA = 1'b0;
            15'b10101110_1010_110: DATA = 1'b0;
            15'b10101110_1010_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 1 Row 11
            15'b10101110_1011_000: DATA = 1'b0;
            15'b10101110_1011_001: DATA = 1'b0;
            15'b10101110_1011_010: DATA = 1'b0;
            15'b10101110_1011_011: DATA = 1'b0;
            15'b10101110_1011_100: DATA = 1'b0;
            15'b10101110_1011_101: DATA = 1'b0;
            15'b10101110_1011_110: DATA = 1'b0;
            15'b10101110_1011_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 1 Row 12
            15'b10101110_1100_000: DATA = 1'b0;
            15'b10101110_1100_001: DATA = 1'b0;
            15'b10101110_1100_010: DATA = 1'b0;
            15'b10101110_1100_011: DATA = 1'b0;
            15'b10101110_1100_100: DATA = 1'b0;
            15'b10101110_1100_101: DATA = 1'b0;
            15'b10101110_1100_110: DATA = 1'b0;
            15'b10101110_1100_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 1 Row 13
            15'b10101110_1101_000: DATA = 1'b0;
            15'b10101110_1101_001: DATA = 1'b0;
            15'b10101110_1101_010: DATA = 1'b0;
            15'b10101110_1101_011: DATA = 1'b0;
            15'b10101110_1101_100: DATA = 1'b0;
            15'b10101110_1101_101: DATA = 1'b0;
            15'b10101110_1101_110: DATA = 1'b0;
            15'b10101110_1101_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 1 Row 14
            15'b10101110_1110_000: DATA = 1'b0;
            15'b10101110_1110_001: DATA = 1'b0;
            15'b10101110_1110_010: DATA = 1'b0;
            15'b10101110_1110_011: DATA = 1'b0;
            15'b10101110_1110_100: DATA = 1'b0;
            15'b10101110_1110_101: DATA = 1'b0;
            15'b10101110_1110_110: DATA = 1'b0;
            15'b10101110_1110_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 1 Row 15
            15'b10101110_1111_000: DATA = 1'b0;
            15'b10101110_1111_001: DATA = 1'b0;
            15'b10101110_1111_010: DATA = 1'b0;
            15'b10101110_1111_011: DATA = 1'b0;
            15'b10101110_1111_100: DATA = 1'b0;
            15'b10101110_1111_101: DATA = 1'b0;
            15'b10101110_1111_110: DATA = 1'b0;
            15'b10101110_1111_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 2 Row 0
            15'b10101111_0000_000: DATA = 1'b0;
            15'b10101111_0000_001: DATA = 1'b0;
            15'b10101111_0000_010: DATA = 1'b0;
            15'b10101111_0000_011: DATA = 1'b0;
            15'b10101111_0000_100: DATA = 1'b0;
            15'b10101111_0000_101: DATA = 1'b0;
            15'b10101111_0000_110: DATA = 1'b0;
            15'b10101111_0000_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 2 Row 1
            15'b10101111_0001_000: DATA = 1'b0;
            15'b10101111_0001_001: DATA = 1'b0;
            15'b10101111_0001_010: DATA = 1'b0;
            15'b10101111_0001_011: DATA = 1'b0;
            15'b10101111_0001_100: DATA = 1'b0;
            15'b10101111_0001_101: DATA = 1'b0;
            15'b10101111_0001_110: DATA = 1'b0;
            15'b10101111_0001_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 2 Row 2
            15'b10101111_0010_000: DATA = 1'b0;
            15'b10101111_0010_001: DATA = 1'b0;
            15'b10101111_0010_010: DATA = 1'b0;
            15'b10101111_0010_011: DATA = 1'b0;
            15'b10101111_0010_100: DATA = 1'b0;
            15'b10101111_0010_101: DATA = 1'b0;
            15'b10101111_0010_110: DATA = 1'b0;
            15'b10101111_0010_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 2 Row 3
            15'b10101111_0011_000: DATA = 1'b0;
            15'b10101111_0011_001: DATA = 1'b0;
            15'b10101111_0011_010: DATA = 1'b0;
            15'b10101111_0011_011: DATA = 1'b0;
            15'b10101111_0011_100: DATA = 1'b0;
            15'b10101111_0011_101: DATA = 1'b0;
            15'b10101111_0011_110: DATA = 1'b0;
            15'b10101111_0011_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 2 Row 4
            15'b10101111_0100_000: DATA = 1'b0;
            15'b10101111_0100_001: DATA = 1'b0;
            15'b10101111_0100_010: DATA = 1'b0;
            15'b10101111_0100_011: DATA = 1'b0;
            15'b10101111_0100_100: DATA = 1'b0;
            15'b10101111_0100_101: DATA = 1'b0;
            15'b10101111_0100_110: DATA = 1'b0;
            15'b10101111_0100_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 2 Row 5
            15'b10101111_0101_000: DATA = 1'b0;
            15'b10101111_0101_001: DATA = 1'b0;
            15'b10101111_0101_010: DATA = 1'b0;
            15'b10101111_0101_011: DATA = 1'b0;
            15'b10101111_0101_100: DATA = 1'b0;
            15'b10101111_0101_101: DATA = 1'b0;
            15'b10101111_0101_110: DATA = 1'b0;
            15'b10101111_0101_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 2 Row 6
            15'b10101111_0110_000: DATA = 1'b0;
            15'b10101111_0110_001: DATA = 1'b0;
            15'b10101111_0110_010: DATA = 1'b0;
            15'b10101111_0110_011: DATA = 1'b0;
            15'b10101111_0110_100: DATA = 1'b0;
            15'b10101111_0110_101: DATA = 1'b0;
            15'b10101111_0110_110: DATA = 1'b0;
            15'b10101111_0110_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 2 Row 7
            15'b10101111_0111_000: DATA = 1'b0;
            15'b10101111_0111_001: DATA = 1'b0;
            15'b10101111_0111_010: DATA = 1'b0;
            15'b10101111_0111_011: DATA = 1'b0;
            15'b10101111_0111_100: DATA = 1'b0;
            15'b10101111_0111_101: DATA = 1'b0;
            15'b10101111_0111_110: DATA = 1'b0;
            15'b10101111_0111_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 2 Row 8
            15'b10101111_1000_000: DATA = 1'b0;
            15'b10101111_1000_001: DATA = 1'b0;
            15'b10101111_1000_010: DATA = 1'b0;
            15'b10101111_1000_011: DATA = 1'b0;
            15'b10101111_1000_100: DATA = 1'b0;
            15'b10101111_1000_101: DATA = 1'b0;
            15'b10101111_1000_110: DATA = 1'b0;
            15'b10101111_1000_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 2 Row 9
            15'b10101111_1001_000: DATA = 1'b0;
            15'b10101111_1001_001: DATA = 1'b0;
            15'b10101111_1001_010: DATA = 1'b0;
            15'b10101111_1001_011: DATA = 1'b0;
            15'b10101111_1001_100: DATA = 1'b0;
            15'b10101111_1001_101: DATA = 1'b0;
            15'b10101111_1001_110: DATA = 1'b0;
            15'b10101111_1001_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 2 Row 10
            15'b10101111_1010_000: DATA = 1'b0;
            15'b10101111_1010_001: DATA = 1'b0;
            15'b10101111_1010_010: DATA = 1'b0;
            15'b10101111_1010_011: DATA = 1'b0;
            15'b10101111_1010_100: DATA = 1'b0;
            15'b10101111_1010_101: DATA = 1'b0;
            15'b10101111_1010_110: DATA = 1'b0;
            15'b10101111_1010_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 2 Row 11
            15'b10101111_1011_000: DATA = 1'b0;
            15'b10101111_1011_001: DATA = 1'b0;
            15'b10101111_1011_010: DATA = 1'b0;
            15'b10101111_1011_011: DATA = 1'b0;
            15'b10101111_1011_100: DATA = 1'b0;
            15'b10101111_1011_101: DATA = 1'b0;
            15'b10101111_1011_110: DATA = 1'b0;
            15'b10101111_1011_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 2 Row 12
            15'b10101111_1100_000: DATA = 1'b0;
            15'b10101111_1100_001: DATA = 1'b0;
            15'b10101111_1100_010: DATA = 1'b0;
            15'b10101111_1100_011: DATA = 1'b0;
            15'b10101111_1100_100: DATA = 1'b0;
            15'b10101111_1100_101: DATA = 1'b0;
            15'b10101111_1100_110: DATA = 1'b0;
            15'b10101111_1100_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 2 Row 13
            15'b10101111_1101_000: DATA = 1'b0;
            15'b10101111_1101_001: DATA = 1'b0;
            15'b10101111_1101_010: DATA = 1'b0;
            15'b10101111_1101_011: DATA = 1'b0;
            15'b10101111_1101_100: DATA = 1'b0;
            15'b10101111_1101_101: DATA = 1'b0;
            15'b10101111_1101_110: DATA = 1'b0;
            15'b10101111_1101_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 2 Row 14
            15'b10101111_1110_000: DATA = 1'b0;
            15'b10101111_1110_001: DATA = 1'b0;
            15'b10101111_1110_010: DATA = 1'b0;
            15'b10101111_1110_011: DATA = 1'b0;
            15'b10101111_1110_100: DATA = 1'b0;
            15'b10101111_1110_101: DATA = 1'b0;
            15'b10101111_1110_110: DATA = 1'b0;
            15'b10101111_1110_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 2 Row 15
            15'b10101111_1111_000: DATA = 1'b0;
            15'b10101111_1111_001: DATA = 1'b0;
            15'b10101111_1111_010: DATA = 1'b0;
            15'b10101111_1111_011: DATA = 1'b0;
            15'b10101111_1111_100: DATA = 1'b0;
            15'b10101111_1111_101: DATA = 1'b0;
            15'b10101111_1111_110: DATA = 1'b0;
            15'b10101111_1111_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 3 Row 0
            15'b10110000_0000_000: DATA = 1'b0;
            15'b10110000_0000_001: DATA = 1'b0;
            15'b10110000_0000_010: DATA = 1'b0;
            15'b10110000_0000_011: DATA = 1'b0;
            15'b10110000_0000_100: DATA = 1'b0;
            15'b10110000_0000_101: DATA = 1'b0;
            15'b10110000_0000_110: DATA = 1'b1;
            15'b10110000_0000_111: DATA = 1'b1;
            // TRIANGLE+ ROW 1 COL 3 Row 1
            15'b10110000_0001_000: DATA = 1'b0;
            15'b10110000_0001_001: DATA = 1'b0;
            15'b10110000_0001_010: DATA = 1'b0;
            15'b10110000_0001_011: DATA = 1'b0;
            15'b10110000_0001_100: DATA = 1'b0;
            15'b10110000_0001_101: DATA = 1'b0;
            15'b10110000_0001_110: DATA = 1'b0;
            15'b10110000_0001_111: DATA = 1'b1;
            // TRIANGLE+ ROW 1 COL 3 Row 2
            15'b10110000_0010_000: DATA = 1'b0;
            15'b10110000_0010_001: DATA = 1'b0;
            15'b10110000_0010_010: DATA = 1'b0;
            15'b10110000_0010_011: DATA = 1'b0;
            15'b10110000_0010_100: DATA = 1'b0;
            15'b10110000_0010_101: DATA = 1'b0;
            15'b10110000_0010_110: DATA = 1'b0;
            15'b10110000_0010_111: DATA = 1'b1;
            // TRIANGLE+ ROW 1 COL 3 Row 3
            15'b10110000_0011_000: DATA = 1'b0;
            15'b10110000_0011_001: DATA = 1'b0;
            15'b10110000_0011_010: DATA = 1'b0;
            15'b10110000_0011_011: DATA = 1'b0;
            15'b10110000_0011_100: DATA = 1'b0;
            15'b10110000_0011_101: DATA = 1'b0;
            15'b10110000_0011_110: DATA = 1'b0;
            15'b10110000_0011_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 3 Row 4
            15'b10110000_0100_000: DATA = 1'b0;
            15'b10110000_0100_001: DATA = 1'b0;
            15'b10110000_0100_010: DATA = 1'b0;
            15'b10110000_0100_011: DATA = 1'b0;
            15'b10110000_0100_100: DATA = 1'b0;
            15'b10110000_0100_101: DATA = 1'b0;
            15'b10110000_0100_110: DATA = 1'b0;
            15'b10110000_0100_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 3 Row 5
            15'b10110000_0101_000: DATA = 1'b0;
            15'b10110000_0101_001: DATA = 1'b0;
            15'b10110000_0101_010: DATA = 1'b0;
            15'b10110000_0101_011: DATA = 1'b0;
            15'b10110000_0101_100: DATA = 1'b0;
            15'b10110000_0101_101: DATA = 1'b0;
            15'b10110000_0101_110: DATA = 1'b0;
            15'b10110000_0101_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 3 Row 6
            15'b10110000_0110_000: DATA = 1'b0;
            15'b10110000_0110_001: DATA = 1'b0;
            15'b10110000_0110_010: DATA = 1'b0;
            15'b10110000_0110_011: DATA = 1'b0;
            15'b10110000_0110_100: DATA = 1'b0;
            15'b10110000_0110_101: DATA = 1'b0;
            15'b10110000_0110_110: DATA = 1'b0;
            15'b10110000_0110_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 3 Row 7
            15'b10110000_0111_000: DATA = 1'b0;
            15'b10110000_0111_001: DATA = 1'b0;
            15'b10110000_0111_010: DATA = 1'b0;
            15'b10110000_0111_011: DATA = 1'b0;
            15'b10110000_0111_100: DATA = 1'b0;
            15'b10110000_0111_101: DATA = 1'b0;
            15'b10110000_0111_110: DATA = 1'b0;
            15'b10110000_0111_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 3 Row 8
            15'b10110000_1000_000: DATA = 1'b0;
            15'b10110000_1000_001: DATA = 1'b0;
            15'b10110000_1000_010: DATA = 1'b0;
            15'b10110000_1000_011: DATA = 1'b0;
            15'b10110000_1000_100: DATA = 1'b0;
            15'b10110000_1000_101: DATA = 1'b0;
            15'b10110000_1000_110: DATA = 1'b0;
            15'b10110000_1000_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 3 Row 9
            15'b10110000_1001_000: DATA = 1'b0;
            15'b10110000_1001_001: DATA = 1'b0;
            15'b10110000_1001_010: DATA = 1'b0;
            15'b10110000_1001_011: DATA = 1'b0;
            15'b10110000_1001_100: DATA = 1'b0;
            15'b10110000_1001_101: DATA = 1'b0;
            15'b10110000_1001_110: DATA = 1'b0;
            15'b10110000_1001_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 3 Row 10
            15'b10110000_1010_000: DATA = 1'b0;
            15'b10110000_1010_001: DATA = 1'b0;
            15'b10110000_1010_010: DATA = 1'b0;
            15'b10110000_1010_011: DATA = 1'b0;
            15'b10110000_1010_100: DATA = 1'b0;
            15'b10110000_1010_101: DATA = 1'b0;
            15'b10110000_1010_110: DATA = 1'b0;
            15'b10110000_1010_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 3 Row 11
            15'b10110000_1011_000: DATA = 1'b0;
            15'b10110000_1011_001: DATA = 1'b0;
            15'b10110000_1011_010: DATA = 1'b0;
            15'b10110000_1011_011: DATA = 1'b0;
            15'b10110000_1011_100: DATA = 1'b0;
            15'b10110000_1011_101: DATA = 1'b0;
            15'b10110000_1011_110: DATA = 1'b0;
            15'b10110000_1011_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 3 Row 12
            15'b10110000_1100_000: DATA = 1'b0;
            15'b10110000_1100_001: DATA = 1'b0;
            15'b10110000_1100_010: DATA = 1'b0;
            15'b10110000_1100_011: DATA = 1'b0;
            15'b10110000_1100_100: DATA = 1'b0;
            15'b10110000_1100_101: DATA = 1'b0;
            15'b10110000_1100_110: DATA = 1'b0;
            15'b10110000_1100_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 3 Row 13
            15'b10110000_1101_000: DATA = 1'b0;
            15'b10110000_1101_001: DATA = 1'b0;
            15'b10110000_1101_010: DATA = 1'b0;
            15'b10110000_1101_011: DATA = 1'b0;
            15'b10110000_1101_100: DATA = 1'b0;
            15'b10110000_1101_101: DATA = 1'b0;
            15'b10110000_1101_110: DATA = 1'b0;
            15'b10110000_1101_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 3 Row 14
            15'b10110000_1110_000: DATA = 1'b0;
            15'b10110000_1110_001: DATA = 1'b0;
            15'b10110000_1110_010: DATA = 1'b0;
            15'b10110000_1110_011: DATA = 1'b0;
            15'b10110000_1110_100: DATA = 1'b0;
            15'b10110000_1110_101: DATA = 1'b0;
            15'b10110000_1110_110: DATA = 1'b0;
            15'b10110000_1110_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 3 Row 15
            15'b10110000_1111_000: DATA = 1'b0;
            15'b10110000_1111_001: DATA = 1'b0;
            15'b10110000_1111_010: DATA = 1'b0;
            15'b10110000_1111_011: DATA = 1'b0;
            15'b10110000_1111_100: DATA = 1'b0;
            15'b10110000_1111_101: DATA = 1'b0;
            15'b10110000_1111_110: DATA = 1'b0;
            15'b10110000_1111_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 4 Row 0
            15'b10110001_0000_000: DATA = 1'b0;
            15'b10110001_0000_001: DATA = 1'b0;
            15'b10110001_0000_010: DATA = 1'b0;
            15'b10110001_0000_011: DATA = 1'b0;
            15'b10110001_0000_100: DATA = 1'b0;
            15'b10110001_0000_101: DATA = 1'b0;
            15'b10110001_0000_110: DATA = 1'b0;
            15'b10110001_0000_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 4 Row 1
            15'b10110001_0001_000: DATA = 1'b0;
            15'b10110001_0001_001: DATA = 1'b0;
            15'b10110001_0001_010: DATA = 1'b0;
            15'b10110001_0001_011: DATA = 1'b0;
            15'b10110001_0001_100: DATA = 1'b0;
            15'b10110001_0001_101: DATA = 1'b0;
            15'b10110001_0001_110: DATA = 1'b0;
            15'b10110001_0001_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 4 Row 2
            15'b10110001_0010_000: DATA = 1'b1;
            15'b10110001_0010_001: DATA = 1'b0;
            15'b10110001_0010_010: DATA = 1'b0;
            15'b10110001_0010_011: DATA = 1'b0;
            15'b10110001_0010_100: DATA = 1'b0;
            15'b10110001_0010_101: DATA = 1'b0;
            15'b10110001_0010_110: DATA = 1'b0;
            15'b10110001_0010_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 4 Row 3
            15'b10110001_0011_000: DATA = 1'b1;
            15'b10110001_0011_001: DATA = 1'b0;
            15'b10110001_0011_010: DATA = 1'b0;
            15'b10110001_0011_011: DATA = 1'b0;
            15'b10110001_0011_100: DATA = 1'b0;
            15'b10110001_0011_101: DATA = 1'b0;
            15'b10110001_0011_110: DATA = 1'b0;
            15'b10110001_0011_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 4 Row 4
            15'b10110001_0100_000: DATA = 1'b1;
            15'b10110001_0100_001: DATA = 1'b1;
            15'b10110001_0100_010: DATA = 1'b0;
            15'b10110001_0100_011: DATA = 1'b0;
            15'b10110001_0100_100: DATA = 1'b0;
            15'b10110001_0100_101: DATA = 1'b0;
            15'b10110001_0100_110: DATA = 1'b0;
            15'b10110001_0100_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 4 Row 5
            15'b10110001_0101_000: DATA = 1'b0;
            15'b10110001_0101_001: DATA = 1'b1;
            15'b10110001_0101_010: DATA = 1'b1;
            15'b10110001_0101_011: DATA = 1'b0;
            15'b10110001_0101_100: DATA = 1'b0;
            15'b10110001_0101_101: DATA = 1'b0;
            15'b10110001_0101_110: DATA = 1'b0;
            15'b10110001_0101_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 4 Row 6
            15'b10110001_0110_000: DATA = 1'b0;
            15'b10110001_0110_001: DATA = 1'b0;
            15'b10110001_0110_010: DATA = 1'b1;
            15'b10110001_0110_011: DATA = 1'b0;
            15'b10110001_0110_100: DATA = 1'b0;
            15'b10110001_0110_101: DATA = 1'b0;
            15'b10110001_0110_110: DATA = 1'b0;
            15'b10110001_0110_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 4 Row 7
            15'b10110001_0111_000: DATA = 1'b0;
            15'b10110001_0111_001: DATA = 1'b0;
            15'b10110001_0111_010: DATA = 1'b1;
            15'b10110001_0111_011: DATA = 1'b1;
            15'b10110001_0111_100: DATA = 1'b0;
            15'b10110001_0111_101: DATA = 1'b0;
            15'b10110001_0111_110: DATA = 1'b0;
            15'b10110001_0111_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 4 Row 8
            15'b10110001_1000_000: DATA = 1'b0;
            15'b10110001_1000_001: DATA = 1'b0;
            15'b10110001_1000_010: DATA = 1'b0;
            15'b10110001_1000_011: DATA = 1'b1;
            15'b10110001_1000_100: DATA = 1'b0;
            15'b10110001_1000_101: DATA = 1'b0;
            15'b10110001_1000_110: DATA = 1'b0;
            15'b10110001_1000_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 4 Row 9
            15'b10110001_1001_000: DATA = 1'b0;
            15'b10110001_1001_001: DATA = 1'b0;
            15'b10110001_1001_010: DATA = 1'b0;
            15'b10110001_1001_011: DATA = 1'b1;
            15'b10110001_1001_100: DATA = 1'b1;
            15'b10110001_1001_101: DATA = 1'b0;
            15'b10110001_1001_110: DATA = 1'b0;
            15'b10110001_1001_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 4 Row 10
            15'b10110001_1010_000: DATA = 1'b0;
            15'b10110001_1010_001: DATA = 1'b0;
            15'b10110001_1010_010: DATA = 1'b0;
            15'b10110001_1010_011: DATA = 1'b0;
            15'b10110001_1010_100: DATA = 1'b1;
            15'b10110001_1010_101: DATA = 1'b1;
            15'b10110001_1010_110: DATA = 1'b0;
            15'b10110001_1010_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 4 Row 11
            15'b10110001_1011_000: DATA = 1'b0;
            15'b10110001_1011_001: DATA = 1'b0;
            15'b10110001_1011_010: DATA = 1'b0;
            15'b10110001_1011_011: DATA = 1'b0;
            15'b10110001_1011_100: DATA = 1'b0;
            15'b10110001_1011_101: DATA = 1'b1;
            15'b10110001_1011_110: DATA = 1'b0;
            15'b10110001_1011_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 4 Row 12
            15'b10110001_1100_000: DATA = 1'b0;
            15'b10110001_1100_001: DATA = 1'b0;
            15'b10110001_1100_010: DATA = 1'b0;
            15'b10110001_1100_011: DATA = 1'b0;
            15'b10110001_1100_100: DATA = 1'b0;
            15'b10110001_1100_101: DATA = 1'b1;
            15'b10110001_1100_110: DATA = 1'b1;
            15'b10110001_1100_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 4 Row 13
            15'b10110001_1101_000: DATA = 1'b0;
            15'b10110001_1101_001: DATA = 1'b0;
            15'b10110001_1101_010: DATA = 1'b0;
            15'b10110001_1101_011: DATA = 1'b0;
            15'b10110001_1101_100: DATA = 1'b0;
            15'b10110001_1101_101: DATA = 1'b0;
            15'b10110001_1101_110: DATA = 1'b1;
            15'b10110001_1101_111: DATA = 1'b0;
            // TRIANGLE+ ROW 1 COL 4 Row 14
            15'b10110001_1110_000: DATA = 1'b0;
            15'b10110001_1110_001: DATA = 1'b0;
            15'b10110001_1110_010: DATA = 1'b0;
            15'b10110001_1110_011: DATA = 1'b0;
            15'b10110001_1110_100: DATA = 1'b0;
            15'b10110001_1110_101: DATA = 1'b0;
            15'b10110001_1110_110: DATA = 1'b1;
            15'b10110001_1110_111: DATA = 1'b1;
            // TRIANGLE+ ROW 1 COL 4 Row 15
            15'b10110001_1111_000: DATA = 1'b0;
            15'b10110001_1111_001: DATA = 1'b0;
            15'b10110001_1111_010: DATA = 1'b0;
            15'b10110001_1111_011: DATA = 1'b0;
            15'b10110001_1111_100: DATA = 1'b0;
            15'b10110001_1111_101: DATA = 1'b0;
            15'b10110001_1111_110: DATA = 1'b0;
            15'b10110001_1111_111: DATA = 1'b1;
            // TRIANGLE- ROW 0 COL 0 Row 0
            15'b10110010_0000_000: DATA = 1'b1;
            15'b10110010_0000_001: DATA = 1'b0;
            15'b10110010_0000_010: DATA = 1'b0;
            15'b10110010_0000_011: DATA = 1'b0;
            15'b10110010_0000_100: DATA = 1'b0;
            15'b10110010_0000_101: DATA = 1'b0;
            15'b10110010_0000_110: DATA = 1'b0;
            15'b10110010_0000_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 0 Row 1
            15'b10110010_0001_000: DATA = 1'b1;
            15'b10110010_0001_001: DATA = 1'b1;
            15'b10110010_0001_010: DATA = 1'b0;
            15'b10110010_0001_011: DATA = 1'b0;
            15'b10110010_0001_100: DATA = 1'b0;
            15'b10110010_0001_101: DATA = 1'b0;
            15'b10110010_0001_110: DATA = 1'b0;
            15'b10110010_0001_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 0 Row 2
            15'b10110010_0010_000: DATA = 1'b0;
            15'b10110010_0010_001: DATA = 1'b1;
            15'b10110010_0010_010: DATA = 1'b0;
            15'b10110010_0010_011: DATA = 1'b0;
            15'b10110010_0010_100: DATA = 1'b0;
            15'b10110010_0010_101: DATA = 1'b0;
            15'b10110010_0010_110: DATA = 1'b0;
            15'b10110010_0010_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 0 Row 3
            15'b10110010_0011_000: DATA = 1'b0;
            15'b10110010_0011_001: DATA = 1'b1;
            15'b10110010_0011_010: DATA = 1'b1;
            15'b10110010_0011_011: DATA = 1'b0;
            15'b10110010_0011_100: DATA = 1'b0;
            15'b10110010_0011_101: DATA = 1'b0;
            15'b10110010_0011_110: DATA = 1'b0;
            15'b10110010_0011_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 0 Row 4
            15'b10110010_0100_000: DATA = 1'b0;
            15'b10110010_0100_001: DATA = 1'b0;
            15'b10110010_0100_010: DATA = 1'b1;
            15'b10110010_0100_011: DATA = 1'b0;
            15'b10110010_0100_100: DATA = 1'b0;
            15'b10110010_0100_101: DATA = 1'b0;
            15'b10110010_0100_110: DATA = 1'b0;
            15'b10110010_0100_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 0 Row 5
            15'b10110010_0101_000: DATA = 1'b0;
            15'b10110010_0101_001: DATA = 1'b0;
            15'b10110010_0101_010: DATA = 1'b1;
            15'b10110010_0101_011: DATA = 1'b1;
            15'b10110010_0101_100: DATA = 1'b0;
            15'b10110010_0101_101: DATA = 1'b0;
            15'b10110010_0101_110: DATA = 1'b0;
            15'b10110010_0101_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 0 Row 6
            15'b10110010_0110_000: DATA = 1'b0;
            15'b10110010_0110_001: DATA = 1'b0;
            15'b10110010_0110_010: DATA = 1'b0;
            15'b10110010_0110_011: DATA = 1'b1;
            15'b10110010_0110_100: DATA = 1'b1;
            15'b10110010_0110_101: DATA = 1'b0;
            15'b10110010_0110_110: DATA = 1'b0;
            15'b10110010_0110_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 0 Row 7
            15'b10110010_0111_000: DATA = 1'b0;
            15'b10110010_0111_001: DATA = 1'b0;
            15'b10110010_0111_010: DATA = 1'b0;
            15'b10110010_0111_011: DATA = 1'b0;
            15'b10110010_0111_100: DATA = 1'b1;
            15'b10110010_0111_101: DATA = 1'b0;
            15'b10110010_0111_110: DATA = 1'b0;
            15'b10110010_0111_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 0 Row 8
            15'b10110010_1000_000: DATA = 1'b0;
            15'b10110010_1000_001: DATA = 1'b0;
            15'b10110010_1000_010: DATA = 1'b0;
            15'b10110010_1000_011: DATA = 1'b0;
            15'b10110010_1000_100: DATA = 1'b1;
            15'b10110010_1000_101: DATA = 1'b1;
            15'b10110010_1000_110: DATA = 1'b0;
            15'b10110010_1000_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 0 Row 9
            15'b10110010_1001_000: DATA = 1'b0;
            15'b10110010_1001_001: DATA = 1'b0;
            15'b10110010_1001_010: DATA = 1'b0;
            15'b10110010_1001_011: DATA = 1'b0;
            15'b10110010_1001_100: DATA = 1'b0;
            15'b10110010_1001_101: DATA = 1'b1;
            15'b10110010_1001_110: DATA = 1'b0;
            15'b10110010_1001_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 0 Row 10
            15'b10110010_1010_000: DATA = 1'b0;
            15'b10110010_1010_001: DATA = 1'b0;
            15'b10110010_1010_010: DATA = 1'b0;
            15'b10110010_1010_011: DATA = 1'b0;
            15'b10110010_1010_100: DATA = 1'b0;
            15'b10110010_1010_101: DATA = 1'b1;
            15'b10110010_1010_110: DATA = 1'b1;
            15'b10110010_1010_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 0 Row 11
            15'b10110010_1011_000: DATA = 1'b0;
            15'b10110010_1011_001: DATA = 1'b0;
            15'b10110010_1011_010: DATA = 1'b0;
            15'b10110010_1011_011: DATA = 1'b0;
            15'b10110010_1011_100: DATA = 1'b0;
            15'b10110010_1011_101: DATA = 1'b0;
            15'b10110010_1011_110: DATA = 1'b1;
            15'b10110010_1011_111: DATA = 1'b1;
            // TRIANGLE- ROW 0 COL 0 Row 12
            15'b10110010_1100_000: DATA = 1'b0;
            15'b10110010_1100_001: DATA = 1'b0;
            15'b10110010_1100_010: DATA = 1'b0;
            15'b10110010_1100_011: DATA = 1'b0;
            15'b10110010_1100_100: DATA = 1'b0;
            15'b10110010_1100_101: DATA = 1'b0;
            15'b10110010_1100_110: DATA = 1'b0;
            15'b10110010_1100_111: DATA = 1'b1;
            // TRIANGLE- ROW 0 COL 0 Row 13
            15'b10110010_1101_000: DATA = 1'b0;
            15'b10110010_1101_001: DATA = 1'b0;
            15'b10110010_1101_010: DATA = 1'b0;
            15'b10110010_1101_011: DATA = 1'b0;
            15'b10110010_1101_100: DATA = 1'b0;
            15'b10110010_1101_101: DATA = 1'b0;
            15'b10110010_1101_110: DATA = 1'b0;
            15'b10110010_1101_111: DATA = 1'b1;
            // TRIANGLE- ROW 0 COL 0 Row 14
            15'b10110010_1110_000: DATA = 1'b0;
            15'b10110010_1110_001: DATA = 1'b0;
            15'b10110010_1110_010: DATA = 1'b0;
            15'b10110010_1110_011: DATA = 1'b0;
            15'b10110010_1110_100: DATA = 1'b0;
            15'b10110010_1110_101: DATA = 1'b0;
            15'b10110010_1110_110: DATA = 1'b0;
            15'b10110010_1110_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 0 Row 15
            15'b10110010_1111_000: DATA = 1'b0;
            15'b10110010_1111_001: DATA = 1'b0;
            15'b10110010_1111_010: DATA = 1'b0;
            15'b10110010_1111_011: DATA = 1'b0;
            15'b10110010_1111_100: DATA = 1'b0;
            15'b10110010_1111_101: DATA = 1'b0;
            15'b10110010_1111_110: DATA = 1'b0;
            15'b10110010_1111_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 1 Row 0
            15'b10110011_0000_000: DATA = 1'b0;
            15'b10110011_0000_001: DATA = 1'b0;
            15'b10110011_0000_010: DATA = 1'b0;
            15'b10110011_0000_011: DATA = 1'b0;
            15'b10110011_0000_100: DATA = 1'b0;
            15'b10110011_0000_101: DATA = 1'b0;
            15'b10110011_0000_110: DATA = 1'b0;
            15'b10110011_0000_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 1 Row 1
            15'b10110011_0001_000: DATA = 1'b0;
            15'b10110011_0001_001: DATA = 1'b0;
            15'b10110011_0001_010: DATA = 1'b0;
            15'b10110011_0001_011: DATA = 1'b0;
            15'b10110011_0001_100: DATA = 1'b0;
            15'b10110011_0001_101: DATA = 1'b0;
            15'b10110011_0001_110: DATA = 1'b0;
            15'b10110011_0001_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 1 Row 2
            15'b10110011_0010_000: DATA = 1'b0;
            15'b10110011_0010_001: DATA = 1'b0;
            15'b10110011_0010_010: DATA = 1'b0;
            15'b10110011_0010_011: DATA = 1'b0;
            15'b10110011_0010_100: DATA = 1'b0;
            15'b10110011_0010_101: DATA = 1'b0;
            15'b10110011_0010_110: DATA = 1'b0;
            15'b10110011_0010_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 1 Row 3
            15'b10110011_0011_000: DATA = 1'b0;
            15'b10110011_0011_001: DATA = 1'b0;
            15'b10110011_0011_010: DATA = 1'b0;
            15'b10110011_0011_011: DATA = 1'b0;
            15'b10110011_0011_100: DATA = 1'b0;
            15'b10110011_0011_101: DATA = 1'b0;
            15'b10110011_0011_110: DATA = 1'b0;
            15'b10110011_0011_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 1 Row 4
            15'b10110011_0100_000: DATA = 1'b0;
            15'b10110011_0100_001: DATA = 1'b0;
            15'b10110011_0100_010: DATA = 1'b0;
            15'b10110011_0100_011: DATA = 1'b0;
            15'b10110011_0100_100: DATA = 1'b0;
            15'b10110011_0100_101: DATA = 1'b0;
            15'b10110011_0100_110: DATA = 1'b0;
            15'b10110011_0100_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 1 Row 5
            15'b10110011_0101_000: DATA = 1'b0;
            15'b10110011_0101_001: DATA = 1'b0;
            15'b10110011_0101_010: DATA = 1'b0;
            15'b10110011_0101_011: DATA = 1'b0;
            15'b10110011_0101_100: DATA = 1'b0;
            15'b10110011_0101_101: DATA = 1'b0;
            15'b10110011_0101_110: DATA = 1'b0;
            15'b10110011_0101_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 1 Row 6
            15'b10110011_0110_000: DATA = 1'b0;
            15'b10110011_0110_001: DATA = 1'b0;
            15'b10110011_0110_010: DATA = 1'b0;
            15'b10110011_0110_011: DATA = 1'b0;
            15'b10110011_0110_100: DATA = 1'b0;
            15'b10110011_0110_101: DATA = 1'b0;
            15'b10110011_0110_110: DATA = 1'b0;
            15'b10110011_0110_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 1 Row 7
            15'b10110011_0111_000: DATA = 1'b0;
            15'b10110011_0111_001: DATA = 1'b0;
            15'b10110011_0111_010: DATA = 1'b0;
            15'b10110011_0111_011: DATA = 1'b0;
            15'b10110011_0111_100: DATA = 1'b0;
            15'b10110011_0111_101: DATA = 1'b0;
            15'b10110011_0111_110: DATA = 1'b0;
            15'b10110011_0111_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 1 Row 8
            15'b10110011_1000_000: DATA = 1'b0;
            15'b10110011_1000_001: DATA = 1'b0;
            15'b10110011_1000_010: DATA = 1'b0;
            15'b10110011_1000_011: DATA = 1'b0;
            15'b10110011_1000_100: DATA = 1'b0;
            15'b10110011_1000_101: DATA = 1'b0;
            15'b10110011_1000_110: DATA = 1'b0;
            15'b10110011_1000_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 1 Row 9
            15'b10110011_1001_000: DATA = 1'b0;
            15'b10110011_1001_001: DATA = 1'b0;
            15'b10110011_1001_010: DATA = 1'b0;
            15'b10110011_1001_011: DATA = 1'b0;
            15'b10110011_1001_100: DATA = 1'b0;
            15'b10110011_1001_101: DATA = 1'b0;
            15'b10110011_1001_110: DATA = 1'b0;
            15'b10110011_1001_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 1 Row 10
            15'b10110011_1010_000: DATA = 1'b0;
            15'b10110011_1010_001: DATA = 1'b0;
            15'b10110011_1010_010: DATA = 1'b0;
            15'b10110011_1010_011: DATA = 1'b0;
            15'b10110011_1010_100: DATA = 1'b0;
            15'b10110011_1010_101: DATA = 1'b0;
            15'b10110011_1010_110: DATA = 1'b0;
            15'b10110011_1010_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 1 Row 11
            15'b10110011_1011_000: DATA = 1'b0;
            15'b10110011_1011_001: DATA = 1'b0;
            15'b10110011_1011_010: DATA = 1'b0;
            15'b10110011_1011_011: DATA = 1'b0;
            15'b10110011_1011_100: DATA = 1'b0;
            15'b10110011_1011_101: DATA = 1'b0;
            15'b10110011_1011_110: DATA = 1'b0;
            15'b10110011_1011_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 1 Row 12
            15'b10110011_1100_000: DATA = 1'b0;
            15'b10110011_1100_001: DATA = 1'b0;
            15'b10110011_1100_010: DATA = 1'b0;
            15'b10110011_1100_011: DATA = 1'b0;
            15'b10110011_1100_100: DATA = 1'b0;
            15'b10110011_1100_101: DATA = 1'b0;
            15'b10110011_1100_110: DATA = 1'b0;
            15'b10110011_1100_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 1 Row 13
            15'b10110011_1101_000: DATA = 1'b1;
            15'b10110011_1101_001: DATA = 1'b0;
            15'b10110011_1101_010: DATA = 1'b0;
            15'b10110011_1101_011: DATA = 1'b0;
            15'b10110011_1101_100: DATA = 1'b0;
            15'b10110011_1101_101: DATA = 1'b0;
            15'b10110011_1101_110: DATA = 1'b0;
            15'b10110011_1101_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 1 Row 14
            15'b10110011_1110_000: DATA = 1'b1;
            15'b10110011_1110_001: DATA = 1'b0;
            15'b10110011_1110_010: DATA = 1'b0;
            15'b10110011_1110_011: DATA = 1'b0;
            15'b10110011_1110_100: DATA = 1'b0;
            15'b10110011_1110_101: DATA = 1'b0;
            15'b10110011_1110_110: DATA = 1'b0;
            15'b10110011_1110_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 1 Row 15
            15'b10110011_1111_000: DATA = 1'b1;
            15'b10110011_1111_001: DATA = 1'b1;
            15'b10110011_1111_010: DATA = 1'b0;
            15'b10110011_1111_011: DATA = 1'b0;
            15'b10110011_1111_100: DATA = 1'b0;
            15'b10110011_1111_101: DATA = 1'b0;
            15'b10110011_1111_110: DATA = 1'b0;
            15'b10110011_1111_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 2 Row 0
            15'b10110100_0000_000: DATA = 1'b0;
            15'b10110100_0000_001: DATA = 1'b0;
            15'b10110100_0000_010: DATA = 1'b0;
            15'b10110100_0000_011: DATA = 1'b0;
            15'b10110100_0000_100: DATA = 1'b0;
            15'b10110100_0000_101: DATA = 1'b0;
            15'b10110100_0000_110: DATA = 1'b0;
            15'b10110100_0000_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 2 Row 1
            15'b10110100_0001_000: DATA = 1'b0;
            15'b10110100_0001_001: DATA = 1'b0;
            15'b10110100_0001_010: DATA = 1'b0;
            15'b10110100_0001_011: DATA = 1'b0;
            15'b10110100_0001_100: DATA = 1'b0;
            15'b10110100_0001_101: DATA = 1'b0;
            15'b10110100_0001_110: DATA = 1'b0;
            15'b10110100_0001_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 2 Row 2
            15'b10110100_0010_000: DATA = 1'b0;
            15'b10110100_0010_001: DATA = 1'b0;
            15'b10110100_0010_010: DATA = 1'b0;
            15'b10110100_0010_011: DATA = 1'b0;
            15'b10110100_0010_100: DATA = 1'b0;
            15'b10110100_0010_101: DATA = 1'b0;
            15'b10110100_0010_110: DATA = 1'b0;
            15'b10110100_0010_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 2 Row 3
            15'b10110100_0011_000: DATA = 1'b0;
            15'b10110100_0011_001: DATA = 1'b0;
            15'b10110100_0011_010: DATA = 1'b0;
            15'b10110100_0011_011: DATA = 1'b0;
            15'b10110100_0011_100: DATA = 1'b0;
            15'b10110100_0011_101: DATA = 1'b0;
            15'b10110100_0011_110: DATA = 1'b0;
            15'b10110100_0011_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 2 Row 4
            15'b10110100_0100_000: DATA = 1'b0;
            15'b10110100_0100_001: DATA = 1'b0;
            15'b10110100_0100_010: DATA = 1'b0;
            15'b10110100_0100_011: DATA = 1'b0;
            15'b10110100_0100_100: DATA = 1'b0;
            15'b10110100_0100_101: DATA = 1'b0;
            15'b10110100_0100_110: DATA = 1'b0;
            15'b10110100_0100_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 2 Row 5
            15'b10110100_0101_000: DATA = 1'b0;
            15'b10110100_0101_001: DATA = 1'b0;
            15'b10110100_0101_010: DATA = 1'b0;
            15'b10110100_0101_011: DATA = 1'b0;
            15'b10110100_0101_100: DATA = 1'b0;
            15'b10110100_0101_101: DATA = 1'b0;
            15'b10110100_0101_110: DATA = 1'b0;
            15'b10110100_0101_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 2 Row 6
            15'b10110100_0110_000: DATA = 1'b0;
            15'b10110100_0110_001: DATA = 1'b0;
            15'b10110100_0110_010: DATA = 1'b0;
            15'b10110100_0110_011: DATA = 1'b0;
            15'b10110100_0110_100: DATA = 1'b0;
            15'b10110100_0110_101: DATA = 1'b0;
            15'b10110100_0110_110: DATA = 1'b0;
            15'b10110100_0110_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 2 Row 7
            15'b10110100_0111_000: DATA = 1'b0;
            15'b10110100_0111_001: DATA = 1'b0;
            15'b10110100_0111_010: DATA = 1'b0;
            15'b10110100_0111_011: DATA = 1'b0;
            15'b10110100_0111_100: DATA = 1'b0;
            15'b10110100_0111_101: DATA = 1'b0;
            15'b10110100_0111_110: DATA = 1'b0;
            15'b10110100_0111_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 2 Row 8
            15'b10110100_1000_000: DATA = 1'b0;
            15'b10110100_1000_001: DATA = 1'b0;
            15'b10110100_1000_010: DATA = 1'b0;
            15'b10110100_1000_011: DATA = 1'b0;
            15'b10110100_1000_100: DATA = 1'b0;
            15'b10110100_1000_101: DATA = 1'b0;
            15'b10110100_1000_110: DATA = 1'b0;
            15'b10110100_1000_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 2 Row 9
            15'b10110100_1001_000: DATA = 1'b0;
            15'b10110100_1001_001: DATA = 1'b0;
            15'b10110100_1001_010: DATA = 1'b0;
            15'b10110100_1001_011: DATA = 1'b0;
            15'b10110100_1001_100: DATA = 1'b0;
            15'b10110100_1001_101: DATA = 1'b0;
            15'b10110100_1001_110: DATA = 1'b0;
            15'b10110100_1001_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 2 Row 10
            15'b10110100_1010_000: DATA = 1'b0;
            15'b10110100_1010_001: DATA = 1'b0;
            15'b10110100_1010_010: DATA = 1'b0;
            15'b10110100_1010_011: DATA = 1'b0;
            15'b10110100_1010_100: DATA = 1'b0;
            15'b10110100_1010_101: DATA = 1'b0;
            15'b10110100_1010_110: DATA = 1'b0;
            15'b10110100_1010_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 2 Row 11
            15'b10110100_1011_000: DATA = 1'b0;
            15'b10110100_1011_001: DATA = 1'b0;
            15'b10110100_1011_010: DATA = 1'b0;
            15'b10110100_1011_011: DATA = 1'b0;
            15'b10110100_1011_100: DATA = 1'b0;
            15'b10110100_1011_101: DATA = 1'b0;
            15'b10110100_1011_110: DATA = 1'b0;
            15'b10110100_1011_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 2 Row 12
            15'b10110100_1100_000: DATA = 1'b0;
            15'b10110100_1100_001: DATA = 1'b0;
            15'b10110100_1100_010: DATA = 1'b0;
            15'b10110100_1100_011: DATA = 1'b0;
            15'b10110100_1100_100: DATA = 1'b0;
            15'b10110100_1100_101: DATA = 1'b0;
            15'b10110100_1100_110: DATA = 1'b0;
            15'b10110100_1100_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 2 Row 13
            15'b10110100_1101_000: DATA = 1'b0;
            15'b10110100_1101_001: DATA = 1'b0;
            15'b10110100_1101_010: DATA = 1'b0;
            15'b10110100_1101_011: DATA = 1'b0;
            15'b10110100_1101_100: DATA = 1'b0;
            15'b10110100_1101_101: DATA = 1'b0;
            15'b10110100_1101_110: DATA = 1'b0;
            15'b10110100_1101_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 2 Row 14
            15'b10110100_1110_000: DATA = 1'b0;
            15'b10110100_1110_001: DATA = 1'b0;
            15'b10110100_1110_010: DATA = 1'b0;
            15'b10110100_1110_011: DATA = 1'b0;
            15'b10110100_1110_100: DATA = 1'b0;
            15'b10110100_1110_101: DATA = 1'b0;
            15'b10110100_1110_110: DATA = 1'b0;
            15'b10110100_1110_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 2 Row 15
            15'b10110100_1111_000: DATA = 1'b0;
            15'b10110100_1111_001: DATA = 1'b0;
            15'b10110100_1111_010: DATA = 1'b0;
            15'b10110100_1111_011: DATA = 1'b0;
            15'b10110100_1111_100: DATA = 1'b0;
            15'b10110100_1111_101: DATA = 1'b0;
            15'b10110100_1111_110: DATA = 1'b0;
            15'b10110100_1111_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 3 Row 0
            15'b10110101_0000_000: DATA = 1'b0;
            15'b10110101_0000_001: DATA = 1'b0;
            15'b10110101_0000_010: DATA = 1'b0;
            15'b10110101_0000_011: DATA = 1'b0;
            15'b10110101_0000_100: DATA = 1'b0;
            15'b10110101_0000_101: DATA = 1'b0;
            15'b10110101_0000_110: DATA = 1'b0;
            15'b10110101_0000_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 3 Row 1
            15'b10110101_0001_000: DATA = 1'b0;
            15'b10110101_0001_001: DATA = 1'b0;
            15'b10110101_0001_010: DATA = 1'b0;
            15'b10110101_0001_011: DATA = 1'b0;
            15'b10110101_0001_100: DATA = 1'b0;
            15'b10110101_0001_101: DATA = 1'b0;
            15'b10110101_0001_110: DATA = 1'b0;
            15'b10110101_0001_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 3 Row 2
            15'b10110101_0010_000: DATA = 1'b0;
            15'b10110101_0010_001: DATA = 1'b0;
            15'b10110101_0010_010: DATA = 1'b0;
            15'b10110101_0010_011: DATA = 1'b0;
            15'b10110101_0010_100: DATA = 1'b0;
            15'b10110101_0010_101: DATA = 1'b0;
            15'b10110101_0010_110: DATA = 1'b0;
            15'b10110101_0010_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 3 Row 3
            15'b10110101_0011_000: DATA = 1'b0;
            15'b10110101_0011_001: DATA = 1'b0;
            15'b10110101_0011_010: DATA = 1'b0;
            15'b10110101_0011_011: DATA = 1'b0;
            15'b10110101_0011_100: DATA = 1'b0;
            15'b10110101_0011_101: DATA = 1'b0;
            15'b10110101_0011_110: DATA = 1'b0;
            15'b10110101_0011_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 3 Row 4
            15'b10110101_0100_000: DATA = 1'b0;
            15'b10110101_0100_001: DATA = 1'b0;
            15'b10110101_0100_010: DATA = 1'b0;
            15'b10110101_0100_011: DATA = 1'b0;
            15'b10110101_0100_100: DATA = 1'b0;
            15'b10110101_0100_101: DATA = 1'b0;
            15'b10110101_0100_110: DATA = 1'b0;
            15'b10110101_0100_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 3 Row 5
            15'b10110101_0101_000: DATA = 1'b0;
            15'b10110101_0101_001: DATA = 1'b0;
            15'b10110101_0101_010: DATA = 1'b0;
            15'b10110101_0101_011: DATA = 1'b0;
            15'b10110101_0101_100: DATA = 1'b0;
            15'b10110101_0101_101: DATA = 1'b0;
            15'b10110101_0101_110: DATA = 1'b0;
            15'b10110101_0101_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 3 Row 6
            15'b10110101_0110_000: DATA = 1'b0;
            15'b10110101_0110_001: DATA = 1'b0;
            15'b10110101_0110_010: DATA = 1'b0;
            15'b10110101_0110_011: DATA = 1'b0;
            15'b10110101_0110_100: DATA = 1'b0;
            15'b10110101_0110_101: DATA = 1'b0;
            15'b10110101_0110_110: DATA = 1'b0;
            15'b10110101_0110_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 3 Row 7
            15'b10110101_0111_000: DATA = 1'b0;
            15'b10110101_0111_001: DATA = 1'b0;
            15'b10110101_0111_010: DATA = 1'b0;
            15'b10110101_0111_011: DATA = 1'b0;
            15'b10110101_0111_100: DATA = 1'b0;
            15'b10110101_0111_101: DATA = 1'b0;
            15'b10110101_0111_110: DATA = 1'b0;
            15'b10110101_0111_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 3 Row 8
            15'b10110101_1000_000: DATA = 1'b0;
            15'b10110101_1000_001: DATA = 1'b0;
            15'b10110101_1000_010: DATA = 1'b0;
            15'b10110101_1000_011: DATA = 1'b0;
            15'b10110101_1000_100: DATA = 1'b0;
            15'b10110101_1000_101: DATA = 1'b0;
            15'b10110101_1000_110: DATA = 1'b0;
            15'b10110101_1000_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 3 Row 9
            15'b10110101_1001_000: DATA = 1'b0;
            15'b10110101_1001_001: DATA = 1'b0;
            15'b10110101_1001_010: DATA = 1'b0;
            15'b10110101_1001_011: DATA = 1'b0;
            15'b10110101_1001_100: DATA = 1'b0;
            15'b10110101_1001_101: DATA = 1'b0;
            15'b10110101_1001_110: DATA = 1'b0;
            15'b10110101_1001_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 3 Row 10
            15'b10110101_1010_000: DATA = 1'b0;
            15'b10110101_1010_001: DATA = 1'b0;
            15'b10110101_1010_010: DATA = 1'b0;
            15'b10110101_1010_011: DATA = 1'b0;
            15'b10110101_1010_100: DATA = 1'b0;
            15'b10110101_1010_101: DATA = 1'b0;
            15'b10110101_1010_110: DATA = 1'b0;
            15'b10110101_1010_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 3 Row 11
            15'b10110101_1011_000: DATA = 1'b0;
            15'b10110101_1011_001: DATA = 1'b0;
            15'b10110101_1011_010: DATA = 1'b0;
            15'b10110101_1011_011: DATA = 1'b0;
            15'b10110101_1011_100: DATA = 1'b0;
            15'b10110101_1011_101: DATA = 1'b0;
            15'b10110101_1011_110: DATA = 1'b0;
            15'b10110101_1011_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 3 Row 12
            15'b10110101_1100_000: DATA = 1'b0;
            15'b10110101_1100_001: DATA = 1'b0;
            15'b10110101_1100_010: DATA = 1'b0;
            15'b10110101_1100_011: DATA = 1'b0;
            15'b10110101_1100_100: DATA = 1'b0;
            15'b10110101_1100_101: DATA = 1'b0;
            15'b10110101_1100_110: DATA = 1'b0;
            15'b10110101_1100_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 3 Row 13
            15'b10110101_1101_000: DATA = 1'b0;
            15'b10110101_1101_001: DATA = 1'b0;
            15'b10110101_1101_010: DATA = 1'b0;
            15'b10110101_1101_011: DATA = 1'b0;
            15'b10110101_1101_100: DATA = 1'b0;
            15'b10110101_1101_101: DATA = 1'b0;
            15'b10110101_1101_110: DATA = 1'b0;
            15'b10110101_1101_111: DATA = 1'b1;
            // TRIANGLE- ROW 0 COL 3 Row 14
            15'b10110101_1110_000: DATA = 1'b0;
            15'b10110101_1110_001: DATA = 1'b0;
            15'b10110101_1110_010: DATA = 1'b0;
            15'b10110101_1110_011: DATA = 1'b0;
            15'b10110101_1110_100: DATA = 1'b0;
            15'b10110101_1110_101: DATA = 1'b0;
            15'b10110101_1110_110: DATA = 1'b0;
            15'b10110101_1110_111: DATA = 1'b1;
            // TRIANGLE- ROW 0 COL 3 Row 15
            15'b10110101_1111_000: DATA = 1'b0;
            15'b10110101_1111_001: DATA = 1'b0;
            15'b10110101_1111_010: DATA = 1'b0;
            15'b10110101_1111_011: DATA = 1'b0;
            15'b10110101_1111_100: DATA = 1'b0;
            15'b10110101_1111_101: DATA = 1'b0;
            15'b10110101_1111_110: DATA = 1'b1;
            15'b10110101_1111_111: DATA = 1'b1;
            // TRIANGLE- ROW 0 COL 4 Row 0
            15'b10110110_0000_000: DATA = 1'b0;
            15'b10110110_0000_001: DATA = 1'b0;
            15'b10110110_0000_010: DATA = 1'b0;
            15'b10110110_0000_011: DATA = 1'b0;
            15'b10110110_0000_100: DATA = 1'b0;
            15'b10110110_0000_101: DATA = 1'b0;
            15'b10110110_0000_110: DATA = 1'b0;
            15'b10110110_0000_111: DATA = 1'b1;
            // TRIANGLE- ROW 0 COL 4 Row 1
            15'b10110110_0001_000: DATA = 1'b0;
            15'b10110110_0001_001: DATA = 1'b0;
            15'b10110110_0001_010: DATA = 1'b0;
            15'b10110110_0001_011: DATA = 1'b0;
            15'b10110110_0001_100: DATA = 1'b0;
            15'b10110110_0001_101: DATA = 1'b0;
            15'b10110110_0001_110: DATA = 1'b1;
            15'b10110110_0001_111: DATA = 1'b1;
            // TRIANGLE- ROW 0 COL 4 Row 2
            15'b10110110_0010_000: DATA = 1'b0;
            15'b10110110_0010_001: DATA = 1'b0;
            15'b10110110_0010_010: DATA = 1'b0;
            15'b10110110_0010_011: DATA = 1'b0;
            15'b10110110_0010_100: DATA = 1'b0;
            15'b10110110_0010_101: DATA = 1'b0;
            15'b10110110_0010_110: DATA = 1'b1;
            15'b10110110_0010_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 4 Row 3
            15'b10110110_0011_000: DATA = 1'b0;
            15'b10110110_0011_001: DATA = 1'b0;
            15'b10110110_0011_010: DATA = 1'b0;
            15'b10110110_0011_011: DATA = 1'b0;
            15'b10110110_0011_100: DATA = 1'b0;
            15'b10110110_0011_101: DATA = 1'b1;
            15'b10110110_0011_110: DATA = 1'b1;
            15'b10110110_0011_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 4 Row 4
            15'b10110110_0100_000: DATA = 1'b0;
            15'b10110110_0100_001: DATA = 1'b0;
            15'b10110110_0100_010: DATA = 1'b0;
            15'b10110110_0100_011: DATA = 1'b0;
            15'b10110110_0100_100: DATA = 1'b0;
            15'b10110110_0100_101: DATA = 1'b1;
            15'b10110110_0100_110: DATA = 1'b0;
            15'b10110110_0100_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 4 Row 5
            15'b10110110_0101_000: DATA = 1'b0;
            15'b10110110_0101_001: DATA = 1'b0;
            15'b10110110_0101_010: DATA = 1'b0;
            15'b10110110_0101_011: DATA = 1'b0;
            15'b10110110_0101_100: DATA = 1'b1;
            15'b10110110_0101_101: DATA = 1'b1;
            15'b10110110_0101_110: DATA = 1'b0;
            15'b10110110_0101_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 4 Row 6
            15'b10110110_0110_000: DATA = 1'b0;
            15'b10110110_0110_001: DATA = 1'b0;
            15'b10110110_0110_010: DATA = 1'b0;
            15'b10110110_0110_011: DATA = 1'b1;
            15'b10110110_0110_100: DATA = 1'b1;
            15'b10110110_0110_101: DATA = 1'b0;
            15'b10110110_0110_110: DATA = 1'b0;
            15'b10110110_0110_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 4 Row 7
            15'b10110110_0111_000: DATA = 1'b0;
            15'b10110110_0111_001: DATA = 1'b0;
            15'b10110110_0111_010: DATA = 1'b0;
            15'b10110110_0111_011: DATA = 1'b1;
            15'b10110110_0111_100: DATA = 1'b0;
            15'b10110110_0111_101: DATA = 1'b0;
            15'b10110110_0111_110: DATA = 1'b0;
            15'b10110110_0111_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 4 Row 8
            15'b10110110_1000_000: DATA = 1'b0;
            15'b10110110_1000_001: DATA = 1'b0;
            15'b10110110_1000_010: DATA = 1'b1;
            15'b10110110_1000_011: DATA = 1'b1;
            15'b10110110_1000_100: DATA = 1'b0;
            15'b10110110_1000_101: DATA = 1'b0;
            15'b10110110_1000_110: DATA = 1'b0;
            15'b10110110_1000_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 4 Row 9
            15'b10110110_1001_000: DATA = 1'b0;
            15'b10110110_1001_001: DATA = 1'b0;
            15'b10110110_1001_010: DATA = 1'b1;
            15'b10110110_1001_011: DATA = 1'b0;
            15'b10110110_1001_100: DATA = 1'b0;
            15'b10110110_1001_101: DATA = 1'b0;
            15'b10110110_1001_110: DATA = 1'b0;
            15'b10110110_1001_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 4 Row 10
            15'b10110110_1010_000: DATA = 1'b0;
            15'b10110110_1010_001: DATA = 1'b1;
            15'b10110110_1010_010: DATA = 1'b1;
            15'b10110110_1010_011: DATA = 1'b0;
            15'b10110110_1010_100: DATA = 1'b0;
            15'b10110110_1010_101: DATA = 1'b0;
            15'b10110110_1010_110: DATA = 1'b0;
            15'b10110110_1010_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 4 Row 11
            15'b10110110_1011_000: DATA = 1'b1;
            15'b10110110_1011_001: DATA = 1'b1;
            15'b10110110_1011_010: DATA = 1'b0;
            15'b10110110_1011_011: DATA = 1'b0;
            15'b10110110_1011_100: DATA = 1'b0;
            15'b10110110_1011_101: DATA = 1'b0;
            15'b10110110_1011_110: DATA = 1'b0;
            15'b10110110_1011_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 4 Row 12
            15'b10110110_1100_000: DATA = 1'b1;
            15'b10110110_1100_001: DATA = 1'b0;
            15'b10110110_1100_010: DATA = 1'b0;
            15'b10110110_1100_011: DATA = 1'b0;
            15'b10110110_1100_100: DATA = 1'b0;
            15'b10110110_1100_101: DATA = 1'b0;
            15'b10110110_1100_110: DATA = 1'b0;
            15'b10110110_1100_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 4 Row 13
            15'b10110110_1101_000: DATA = 1'b1;
            15'b10110110_1101_001: DATA = 1'b0;
            15'b10110110_1101_010: DATA = 1'b0;
            15'b10110110_1101_011: DATA = 1'b0;
            15'b10110110_1101_100: DATA = 1'b0;
            15'b10110110_1101_101: DATA = 1'b0;
            15'b10110110_1101_110: DATA = 1'b0;
            15'b10110110_1101_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 4 Row 14
            15'b10110110_1110_000: DATA = 1'b0;
            15'b10110110_1110_001: DATA = 1'b0;
            15'b10110110_1110_010: DATA = 1'b0;
            15'b10110110_1110_011: DATA = 1'b0;
            15'b10110110_1110_100: DATA = 1'b0;
            15'b10110110_1110_101: DATA = 1'b0;
            15'b10110110_1110_110: DATA = 1'b0;
            15'b10110110_1110_111: DATA = 1'b0;
            // TRIANGLE- ROW 0 COL 4 Row 15
            15'b10110110_1111_000: DATA = 1'b0;
            15'b10110110_1111_001: DATA = 1'b0;
            15'b10110110_1111_010: DATA = 1'b0;
            15'b10110110_1111_011: DATA = 1'b0;
            15'b10110110_1111_100: DATA = 1'b0;
            15'b10110110_1111_101: DATA = 1'b0;
            15'b10110110_1111_110: DATA = 1'b0;
            15'b10110110_1111_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 0 Row 0
            15'b10110111_0000_000: DATA = 1'b0;
            15'b10110111_0000_001: DATA = 1'b0;
            15'b10110111_0000_010: DATA = 1'b0;
            15'b10110111_0000_011: DATA = 1'b0;
            15'b10110111_0000_100: DATA = 1'b0;
            15'b10110111_0000_101: DATA = 1'b0;
            15'b10110111_0000_110: DATA = 1'b0;
            15'b10110111_0000_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 0 Row 1
            15'b10110111_0001_000: DATA = 1'b0;
            15'b10110111_0001_001: DATA = 1'b0;
            15'b10110111_0001_010: DATA = 1'b0;
            15'b10110111_0001_011: DATA = 1'b0;
            15'b10110111_0001_100: DATA = 1'b0;
            15'b10110111_0001_101: DATA = 1'b0;
            15'b10110111_0001_110: DATA = 1'b0;
            15'b10110111_0001_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 0 Row 2
            15'b10110111_0010_000: DATA = 1'b0;
            15'b10110111_0010_001: DATA = 1'b0;
            15'b10110111_0010_010: DATA = 1'b0;
            15'b10110111_0010_011: DATA = 1'b0;
            15'b10110111_0010_100: DATA = 1'b0;
            15'b10110111_0010_101: DATA = 1'b0;
            15'b10110111_0010_110: DATA = 1'b0;
            15'b10110111_0010_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 0 Row 3
            15'b10110111_0011_000: DATA = 1'b0;
            15'b10110111_0011_001: DATA = 1'b0;
            15'b10110111_0011_010: DATA = 1'b0;
            15'b10110111_0011_011: DATA = 1'b0;
            15'b10110111_0011_100: DATA = 1'b0;
            15'b10110111_0011_101: DATA = 1'b0;
            15'b10110111_0011_110: DATA = 1'b0;
            15'b10110111_0011_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 0 Row 4
            15'b10110111_0100_000: DATA = 1'b0;
            15'b10110111_0100_001: DATA = 1'b0;
            15'b10110111_0100_010: DATA = 1'b0;
            15'b10110111_0100_011: DATA = 1'b0;
            15'b10110111_0100_100: DATA = 1'b0;
            15'b10110111_0100_101: DATA = 1'b0;
            15'b10110111_0100_110: DATA = 1'b0;
            15'b10110111_0100_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 0 Row 5
            15'b10110111_0101_000: DATA = 1'b0;
            15'b10110111_0101_001: DATA = 1'b0;
            15'b10110111_0101_010: DATA = 1'b0;
            15'b10110111_0101_011: DATA = 1'b0;
            15'b10110111_0101_100: DATA = 1'b0;
            15'b10110111_0101_101: DATA = 1'b0;
            15'b10110111_0101_110: DATA = 1'b0;
            15'b10110111_0101_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 0 Row 6
            15'b10110111_0110_000: DATA = 1'b0;
            15'b10110111_0110_001: DATA = 1'b0;
            15'b10110111_0110_010: DATA = 1'b0;
            15'b10110111_0110_011: DATA = 1'b0;
            15'b10110111_0110_100: DATA = 1'b0;
            15'b10110111_0110_101: DATA = 1'b0;
            15'b10110111_0110_110: DATA = 1'b0;
            15'b10110111_0110_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 0 Row 7
            15'b10110111_0111_000: DATA = 1'b0;
            15'b10110111_0111_001: DATA = 1'b0;
            15'b10110111_0111_010: DATA = 1'b0;
            15'b10110111_0111_011: DATA = 1'b0;
            15'b10110111_0111_100: DATA = 1'b0;
            15'b10110111_0111_101: DATA = 1'b0;
            15'b10110111_0111_110: DATA = 1'b0;
            15'b10110111_0111_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 0 Row 8
            15'b10110111_1000_000: DATA = 1'b0;
            15'b10110111_1000_001: DATA = 1'b0;
            15'b10110111_1000_010: DATA = 1'b0;
            15'b10110111_1000_011: DATA = 1'b0;
            15'b10110111_1000_100: DATA = 1'b0;
            15'b10110111_1000_101: DATA = 1'b0;
            15'b10110111_1000_110: DATA = 1'b0;
            15'b10110111_1000_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 0 Row 9
            15'b10110111_1001_000: DATA = 1'b0;
            15'b10110111_1001_001: DATA = 1'b0;
            15'b10110111_1001_010: DATA = 1'b0;
            15'b10110111_1001_011: DATA = 1'b0;
            15'b10110111_1001_100: DATA = 1'b0;
            15'b10110111_1001_101: DATA = 1'b0;
            15'b10110111_1001_110: DATA = 1'b0;
            15'b10110111_1001_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 0 Row 10
            15'b10110111_1010_000: DATA = 1'b0;
            15'b10110111_1010_001: DATA = 1'b0;
            15'b10110111_1010_010: DATA = 1'b0;
            15'b10110111_1010_011: DATA = 1'b0;
            15'b10110111_1010_100: DATA = 1'b0;
            15'b10110111_1010_101: DATA = 1'b0;
            15'b10110111_1010_110: DATA = 1'b0;
            15'b10110111_1010_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 0 Row 11
            15'b10110111_1011_000: DATA = 1'b0;
            15'b10110111_1011_001: DATA = 1'b0;
            15'b10110111_1011_010: DATA = 1'b0;
            15'b10110111_1011_011: DATA = 1'b0;
            15'b10110111_1011_100: DATA = 1'b0;
            15'b10110111_1011_101: DATA = 1'b0;
            15'b10110111_1011_110: DATA = 1'b0;
            15'b10110111_1011_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 0 Row 12
            15'b10110111_1100_000: DATA = 1'b0;
            15'b10110111_1100_001: DATA = 1'b0;
            15'b10110111_1100_010: DATA = 1'b0;
            15'b10110111_1100_011: DATA = 1'b0;
            15'b10110111_1100_100: DATA = 1'b0;
            15'b10110111_1100_101: DATA = 1'b0;
            15'b10110111_1100_110: DATA = 1'b0;
            15'b10110111_1100_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 0 Row 13
            15'b10110111_1101_000: DATA = 1'b0;
            15'b10110111_1101_001: DATA = 1'b0;
            15'b10110111_1101_010: DATA = 1'b0;
            15'b10110111_1101_011: DATA = 1'b0;
            15'b10110111_1101_100: DATA = 1'b0;
            15'b10110111_1101_101: DATA = 1'b0;
            15'b10110111_1101_110: DATA = 1'b0;
            15'b10110111_1101_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 0 Row 14
            15'b10110111_1110_000: DATA = 1'b0;
            15'b10110111_1110_001: DATA = 1'b0;
            15'b10110111_1110_010: DATA = 1'b0;
            15'b10110111_1110_011: DATA = 1'b0;
            15'b10110111_1110_100: DATA = 1'b0;
            15'b10110111_1110_101: DATA = 1'b0;
            15'b10110111_1110_110: DATA = 1'b0;
            15'b10110111_1110_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 0 Row 15
            15'b10110111_1111_000: DATA = 1'b0;
            15'b10110111_1111_001: DATA = 1'b0;
            15'b10110111_1111_010: DATA = 1'b0;
            15'b10110111_1111_011: DATA = 1'b0;
            15'b10110111_1111_100: DATA = 1'b0;
            15'b10110111_1111_101: DATA = 1'b0;
            15'b10110111_1111_110: DATA = 1'b0;
            15'b10110111_1111_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 1 Row 0
            15'b10111000_0000_000: DATA = 1'b0;
            15'b10111000_0000_001: DATA = 1'b1;
            15'b10111000_0000_010: DATA = 1'b1;
            15'b10111000_0000_011: DATA = 1'b0;
            15'b10111000_0000_100: DATA = 1'b0;
            15'b10111000_0000_101: DATA = 1'b0;
            15'b10111000_0000_110: DATA = 1'b0;
            15'b10111000_0000_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 1 Row 1
            15'b10111000_0001_000: DATA = 1'b0;
            15'b10111000_0001_001: DATA = 1'b0;
            15'b10111000_0001_010: DATA = 1'b1;
            15'b10111000_0001_011: DATA = 1'b0;
            15'b10111000_0001_100: DATA = 1'b0;
            15'b10111000_0001_101: DATA = 1'b0;
            15'b10111000_0001_110: DATA = 1'b0;
            15'b10111000_0001_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 1 Row 2
            15'b10111000_0010_000: DATA = 1'b0;
            15'b10111000_0010_001: DATA = 1'b0;
            15'b10111000_0010_010: DATA = 1'b1;
            15'b10111000_0010_011: DATA = 1'b1;
            15'b10111000_0010_100: DATA = 1'b0;
            15'b10111000_0010_101: DATA = 1'b0;
            15'b10111000_0010_110: DATA = 1'b0;
            15'b10111000_0010_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 1 Row 3
            15'b10111000_0011_000: DATA = 1'b0;
            15'b10111000_0011_001: DATA = 1'b0;
            15'b10111000_0011_010: DATA = 1'b0;
            15'b10111000_0011_011: DATA = 1'b1;
            15'b10111000_0011_100: DATA = 1'b0;
            15'b10111000_0011_101: DATA = 1'b0;
            15'b10111000_0011_110: DATA = 1'b0;
            15'b10111000_0011_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 1 Row 4
            15'b10111000_0100_000: DATA = 1'b0;
            15'b10111000_0100_001: DATA = 1'b0;
            15'b10111000_0100_010: DATA = 1'b0;
            15'b10111000_0100_011: DATA = 1'b1;
            15'b10111000_0100_100: DATA = 1'b1;
            15'b10111000_0100_101: DATA = 1'b0;
            15'b10111000_0100_110: DATA = 1'b0;
            15'b10111000_0100_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 1 Row 5
            15'b10111000_0101_000: DATA = 1'b0;
            15'b10111000_0101_001: DATA = 1'b0;
            15'b10111000_0101_010: DATA = 1'b0;
            15'b10111000_0101_011: DATA = 1'b0;
            15'b10111000_0101_100: DATA = 1'b1;
            15'b10111000_0101_101: DATA = 1'b1;
            15'b10111000_0101_110: DATA = 1'b0;
            15'b10111000_0101_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 1 Row 6
            15'b10111000_0110_000: DATA = 1'b0;
            15'b10111000_0110_001: DATA = 1'b0;
            15'b10111000_0110_010: DATA = 1'b0;
            15'b10111000_0110_011: DATA = 1'b0;
            15'b10111000_0110_100: DATA = 1'b0;
            15'b10111000_0110_101: DATA = 1'b1;
            15'b10111000_0110_110: DATA = 1'b0;
            15'b10111000_0110_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 1 Row 7
            15'b10111000_0111_000: DATA = 1'b0;
            15'b10111000_0111_001: DATA = 1'b0;
            15'b10111000_0111_010: DATA = 1'b0;
            15'b10111000_0111_011: DATA = 1'b0;
            15'b10111000_0111_100: DATA = 1'b0;
            15'b10111000_0111_101: DATA = 1'b1;
            15'b10111000_0111_110: DATA = 1'b1;
            15'b10111000_0111_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 1 Row 8
            15'b10111000_1000_000: DATA = 1'b0;
            15'b10111000_1000_001: DATA = 1'b0;
            15'b10111000_1000_010: DATA = 1'b0;
            15'b10111000_1000_011: DATA = 1'b0;
            15'b10111000_1000_100: DATA = 1'b0;
            15'b10111000_1000_101: DATA = 1'b0;
            15'b10111000_1000_110: DATA = 1'b1;
            15'b10111000_1000_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 1 Row 9
            15'b10111000_1001_000: DATA = 1'b0;
            15'b10111000_1001_001: DATA = 1'b0;
            15'b10111000_1001_010: DATA = 1'b0;
            15'b10111000_1001_011: DATA = 1'b0;
            15'b10111000_1001_100: DATA = 1'b0;
            15'b10111000_1001_101: DATA = 1'b0;
            15'b10111000_1001_110: DATA = 1'b1;
            15'b10111000_1001_111: DATA = 1'b1;
            // TRIANGLE- ROW 1 COL 1 Row 10
            15'b10111000_1010_000: DATA = 1'b0;
            15'b10111000_1010_001: DATA = 1'b0;
            15'b10111000_1010_010: DATA = 1'b0;
            15'b10111000_1010_011: DATA = 1'b0;
            15'b10111000_1010_100: DATA = 1'b0;
            15'b10111000_1010_101: DATA = 1'b0;
            15'b10111000_1010_110: DATA = 1'b0;
            15'b10111000_1010_111: DATA = 1'b1;
            // TRIANGLE- ROW 1 COL 1 Row 11
            15'b10111000_1011_000: DATA = 1'b0;
            15'b10111000_1011_001: DATA = 1'b0;
            15'b10111000_1011_010: DATA = 1'b0;
            15'b10111000_1011_011: DATA = 1'b0;
            15'b10111000_1011_100: DATA = 1'b0;
            15'b10111000_1011_101: DATA = 1'b0;
            15'b10111000_1011_110: DATA = 1'b0;
            15'b10111000_1011_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 1 Row 12
            15'b10111000_1100_000: DATA = 1'b0;
            15'b10111000_1100_001: DATA = 1'b0;
            15'b10111000_1100_010: DATA = 1'b0;
            15'b10111000_1100_011: DATA = 1'b0;
            15'b10111000_1100_100: DATA = 1'b0;
            15'b10111000_1100_101: DATA = 1'b0;
            15'b10111000_1100_110: DATA = 1'b0;
            15'b10111000_1100_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 1 Row 13
            15'b10111000_1101_000: DATA = 1'b0;
            15'b10111000_1101_001: DATA = 1'b0;
            15'b10111000_1101_010: DATA = 1'b0;
            15'b10111000_1101_011: DATA = 1'b0;
            15'b10111000_1101_100: DATA = 1'b0;
            15'b10111000_1101_101: DATA = 1'b0;
            15'b10111000_1101_110: DATA = 1'b0;
            15'b10111000_1101_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 1 Row 14
            15'b10111000_1110_000: DATA = 1'b0;
            15'b10111000_1110_001: DATA = 1'b0;
            15'b10111000_1110_010: DATA = 1'b0;
            15'b10111000_1110_011: DATA = 1'b0;
            15'b10111000_1110_100: DATA = 1'b0;
            15'b10111000_1110_101: DATA = 1'b0;
            15'b10111000_1110_110: DATA = 1'b0;
            15'b10111000_1110_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 1 Row 15
            15'b10111000_1111_000: DATA = 1'b0;
            15'b10111000_1111_001: DATA = 1'b0;
            15'b10111000_1111_010: DATA = 1'b0;
            15'b10111000_1111_011: DATA = 1'b0;
            15'b10111000_1111_100: DATA = 1'b0;
            15'b10111000_1111_101: DATA = 1'b0;
            15'b10111000_1111_110: DATA = 1'b0;
            15'b10111000_1111_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 2 Row 0
            15'b10111001_0000_000: DATA = 1'b0;
            15'b10111001_0000_001: DATA = 1'b0;
            15'b10111001_0000_010: DATA = 1'b0;
            15'b10111001_0000_011: DATA = 1'b0;
            15'b10111001_0000_100: DATA = 1'b0;
            15'b10111001_0000_101: DATA = 1'b0;
            15'b10111001_0000_110: DATA = 1'b0;
            15'b10111001_0000_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 2 Row 1
            15'b10111001_0001_000: DATA = 1'b0;
            15'b10111001_0001_001: DATA = 1'b0;
            15'b10111001_0001_010: DATA = 1'b0;
            15'b10111001_0001_011: DATA = 1'b0;
            15'b10111001_0001_100: DATA = 1'b0;
            15'b10111001_0001_101: DATA = 1'b0;
            15'b10111001_0001_110: DATA = 1'b0;
            15'b10111001_0001_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 2 Row 2
            15'b10111001_0010_000: DATA = 1'b0;
            15'b10111001_0010_001: DATA = 1'b0;
            15'b10111001_0010_010: DATA = 1'b0;
            15'b10111001_0010_011: DATA = 1'b0;
            15'b10111001_0010_100: DATA = 1'b0;
            15'b10111001_0010_101: DATA = 1'b0;
            15'b10111001_0010_110: DATA = 1'b0;
            15'b10111001_0010_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 2 Row 3
            15'b10111001_0011_000: DATA = 1'b0;
            15'b10111001_0011_001: DATA = 1'b0;
            15'b10111001_0011_010: DATA = 1'b0;
            15'b10111001_0011_011: DATA = 1'b0;
            15'b10111001_0011_100: DATA = 1'b0;
            15'b10111001_0011_101: DATA = 1'b0;
            15'b10111001_0011_110: DATA = 1'b0;
            15'b10111001_0011_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 2 Row 4
            15'b10111001_0100_000: DATA = 1'b0;
            15'b10111001_0100_001: DATA = 1'b0;
            15'b10111001_0100_010: DATA = 1'b0;
            15'b10111001_0100_011: DATA = 1'b0;
            15'b10111001_0100_100: DATA = 1'b0;
            15'b10111001_0100_101: DATA = 1'b0;
            15'b10111001_0100_110: DATA = 1'b0;
            15'b10111001_0100_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 2 Row 5
            15'b10111001_0101_000: DATA = 1'b0;
            15'b10111001_0101_001: DATA = 1'b0;
            15'b10111001_0101_010: DATA = 1'b0;
            15'b10111001_0101_011: DATA = 1'b0;
            15'b10111001_0101_100: DATA = 1'b0;
            15'b10111001_0101_101: DATA = 1'b0;
            15'b10111001_0101_110: DATA = 1'b0;
            15'b10111001_0101_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 2 Row 6
            15'b10111001_0110_000: DATA = 1'b0;
            15'b10111001_0110_001: DATA = 1'b0;
            15'b10111001_0110_010: DATA = 1'b0;
            15'b10111001_0110_011: DATA = 1'b0;
            15'b10111001_0110_100: DATA = 1'b0;
            15'b10111001_0110_101: DATA = 1'b0;
            15'b10111001_0110_110: DATA = 1'b0;
            15'b10111001_0110_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 2 Row 7
            15'b10111001_0111_000: DATA = 1'b0;
            15'b10111001_0111_001: DATA = 1'b0;
            15'b10111001_0111_010: DATA = 1'b0;
            15'b10111001_0111_011: DATA = 1'b0;
            15'b10111001_0111_100: DATA = 1'b0;
            15'b10111001_0111_101: DATA = 1'b0;
            15'b10111001_0111_110: DATA = 1'b0;
            15'b10111001_0111_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 2 Row 8
            15'b10111001_1000_000: DATA = 1'b0;
            15'b10111001_1000_001: DATA = 1'b0;
            15'b10111001_1000_010: DATA = 1'b0;
            15'b10111001_1000_011: DATA = 1'b0;
            15'b10111001_1000_100: DATA = 1'b0;
            15'b10111001_1000_101: DATA = 1'b0;
            15'b10111001_1000_110: DATA = 1'b0;
            15'b10111001_1000_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 2 Row 9
            15'b10111001_1001_000: DATA = 1'b0;
            15'b10111001_1001_001: DATA = 1'b0;
            15'b10111001_1001_010: DATA = 1'b0;
            15'b10111001_1001_011: DATA = 1'b0;
            15'b10111001_1001_100: DATA = 1'b0;
            15'b10111001_1001_101: DATA = 1'b0;
            15'b10111001_1001_110: DATA = 1'b0;
            15'b10111001_1001_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 2 Row 10
            15'b10111001_1010_000: DATA = 1'b1;
            15'b10111001_1010_001: DATA = 1'b0;
            15'b10111001_1010_010: DATA = 1'b0;
            15'b10111001_1010_011: DATA = 1'b0;
            15'b10111001_1010_100: DATA = 1'b0;
            15'b10111001_1010_101: DATA = 1'b0;
            15'b10111001_1010_110: DATA = 1'b0;
            15'b10111001_1010_111: DATA = 1'b1;
            // TRIANGLE- ROW 1 COL 2 Row 11
            15'b10111001_1011_000: DATA = 1'b1;
            15'b10111001_1011_001: DATA = 1'b0;
            15'b10111001_1011_010: DATA = 1'b0;
            15'b10111001_1011_011: DATA = 1'b0;
            15'b10111001_1011_100: DATA = 1'b0;
            15'b10111001_1011_101: DATA = 1'b0;
            15'b10111001_1011_110: DATA = 1'b0;
            15'b10111001_1011_111: DATA = 1'b1;
            // TRIANGLE- ROW 1 COL 2 Row 12
            15'b10111001_1100_000: DATA = 1'b1;
            15'b10111001_1100_001: DATA = 1'b1;
            15'b10111001_1100_010: DATA = 1'b0;
            15'b10111001_1100_011: DATA = 1'b0;
            15'b10111001_1100_100: DATA = 1'b0;
            15'b10111001_1100_101: DATA = 1'b0;
            15'b10111001_1100_110: DATA = 1'b1;
            15'b10111001_1100_111: DATA = 1'b1;
            // TRIANGLE- ROW 1 COL 2 Row 13
            15'b10111001_1101_000: DATA = 1'b0;
            15'b10111001_1101_001: DATA = 1'b1;
            15'b10111001_1101_010: DATA = 1'b0;
            15'b10111001_1101_011: DATA = 1'b0;
            15'b10111001_1101_100: DATA = 1'b0;
            15'b10111001_1101_101: DATA = 1'b0;
            15'b10111001_1101_110: DATA = 1'b1;
            15'b10111001_1101_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 2 Row 14
            15'b10111001_1110_000: DATA = 1'b0;
            15'b10111001_1110_001: DATA = 1'b1;
            15'b10111001_1110_010: DATA = 1'b1;
            15'b10111001_1110_011: DATA = 1'b0;
            15'b10111001_1110_100: DATA = 1'b0;
            15'b10111001_1110_101: DATA = 1'b1;
            15'b10111001_1110_110: DATA = 1'b1;
            15'b10111001_1110_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 2 Row 15
            15'b10111001_1111_000: DATA = 1'b0;
            15'b10111001_1111_001: DATA = 1'b0;
            15'b10111001_1111_010: DATA = 1'b0;
            15'b10111001_1111_011: DATA = 1'b1;
            15'b10111001_1111_100: DATA = 1'b1;
            15'b10111001_1111_101: DATA = 1'b0;
            15'b10111001_1111_110: DATA = 1'b0;
            15'b10111001_1111_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 3 Row 0
            15'b10111010_0000_000: DATA = 1'b0;
            15'b10111010_0000_001: DATA = 1'b0;
            15'b10111010_0000_010: DATA = 1'b0;
            15'b10111010_0000_011: DATA = 1'b0;
            15'b10111010_0000_100: DATA = 1'b0;
            15'b10111010_0000_101: DATA = 1'b1;
            15'b10111010_0000_110: DATA = 1'b1;
            15'b10111010_0000_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 3 Row 1
            15'b10111010_0001_000: DATA = 1'b0;
            15'b10111010_0001_001: DATA = 1'b0;
            15'b10111010_0001_010: DATA = 1'b0;
            15'b10111010_0001_011: DATA = 1'b0;
            15'b10111010_0001_100: DATA = 1'b0;
            15'b10111010_0001_101: DATA = 1'b1;
            15'b10111010_0001_110: DATA = 1'b0;
            15'b10111010_0001_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 3 Row 2
            15'b10111010_0010_000: DATA = 1'b0;
            15'b10111010_0010_001: DATA = 1'b0;
            15'b10111010_0010_010: DATA = 1'b0;
            15'b10111010_0010_011: DATA = 1'b0;
            15'b10111010_0010_100: DATA = 1'b1;
            15'b10111010_0010_101: DATA = 1'b1;
            15'b10111010_0010_110: DATA = 1'b0;
            15'b10111010_0010_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 3 Row 3
            15'b10111010_0011_000: DATA = 1'b0;
            15'b10111010_0011_001: DATA = 1'b0;
            15'b10111010_0011_010: DATA = 1'b0;
            15'b10111010_0011_011: DATA = 1'b0;
            15'b10111010_0011_100: DATA = 1'b1;
            15'b10111010_0011_101: DATA = 1'b0;
            15'b10111010_0011_110: DATA = 1'b0;
            15'b10111010_0011_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 3 Row 4
            15'b10111010_0100_000: DATA = 1'b0;
            15'b10111010_0100_001: DATA = 1'b0;
            15'b10111010_0100_010: DATA = 1'b0;
            15'b10111010_0100_011: DATA = 1'b1;
            15'b10111010_0100_100: DATA = 1'b1;
            15'b10111010_0100_101: DATA = 1'b0;
            15'b10111010_0100_110: DATA = 1'b0;
            15'b10111010_0100_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 3 Row 5
            15'b10111010_0101_000: DATA = 1'b0;
            15'b10111010_0101_001: DATA = 1'b0;
            15'b10111010_0101_010: DATA = 1'b1;
            15'b10111010_0101_011: DATA = 1'b1;
            15'b10111010_0101_100: DATA = 1'b0;
            15'b10111010_0101_101: DATA = 1'b0;
            15'b10111010_0101_110: DATA = 1'b0;
            15'b10111010_0101_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 3 Row 6
            15'b10111010_0110_000: DATA = 1'b0;
            15'b10111010_0110_001: DATA = 1'b0;
            15'b10111010_0110_010: DATA = 1'b1;
            15'b10111010_0110_011: DATA = 1'b0;
            15'b10111010_0110_100: DATA = 1'b0;
            15'b10111010_0110_101: DATA = 1'b0;
            15'b10111010_0110_110: DATA = 1'b0;
            15'b10111010_0110_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 3 Row 7
            15'b10111010_0111_000: DATA = 1'b0;
            15'b10111010_0111_001: DATA = 1'b1;
            15'b10111010_0111_010: DATA = 1'b1;
            15'b10111010_0111_011: DATA = 1'b0;
            15'b10111010_0111_100: DATA = 1'b0;
            15'b10111010_0111_101: DATA = 1'b0;
            15'b10111010_0111_110: DATA = 1'b0;
            15'b10111010_0111_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 3 Row 8
            15'b10111010_1000_000: DATA = 1'b0;
            15'b10111010_1000_001: DATA = 1'b1;
            15'b10111010_1000_010: DATA = 1'b0;
            15'b10111010_1000_011: DATA = 1'b0;
            15'b10111010_1000_100: DATA = 1'b0;
            15'b10111010_1000_101: DATA = 1'b0;
            15'b10111010_1000_110: DATA = 1'b0;
            15'b10111010_1000_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 3 Row 9
            15'b10111010_1001_000: DATA = 1'b1;
            15'b10111010_1001_001: DATA = 1'b1;
            15'b10111010_1001_010: DATA = 1'b0;
            15'b10111010_1001_011: DATA = 1'b0;
            15'b10111010_1001_100: DATA = 1'b0;
            15'b10111010_1001_101: DATA = 1'b0;
            15'b10111010_1001_110: DATA = 1'b0;
            15'b10111010_1001_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 3 Row 10
            15'b10111010_1010_000: DATA = 1'b1;
            15'b10111010_1010_001: DATA = 1'b0;
            15'b10111010_1010_010: DATA = 1'b0;
            15'b10111010_1010_011: DATA = 1'b0;
            15'b10111010_1010_100: DATA = 1'b0;
            15'b10111010_1010_101: DATA = 1'b0;
            15'b10111010_1010_110: DATA = 1'b0;
            15'b10111010_1010_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 3 Row 11
            15'b10111010_1011_000: DATA = 1'b0;
            15'b10111010_1011_001: DATA = 1'b0;
            15'b10111010_1011_010: DATA = 1'b0;
            15'b10111010_1011_011: DATA = 1'b0;
            15'b10111010_1011_100: DATA = 1'b0;
            15'b10111010_1011_101: DATA = 1'b0;
            15'b10111010_1011_110: DATA = 1'b0;
            15'b10111010_1011_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 3 Row 12
            15'b10111010_1100_000: DATA = 1'b0;
            15'b10111010_1100_001: DATA = 1'b0;
            15'b10111010_1100_010: DATA = 1'b0;
            15'b10111010_1100_011: DATA = 1'b0;
            15'b10111010_1100_100: DATA = 1'b0;
            15'b10111010_1100_101: DATA = 1'b0;
            15'b10111010_1100_110: DATA = 1'b0;
            15'b10111010_1100_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 3 Row 13
            15'b10111010_1101_000: DATA = 1'b0;
            15'b10111010_1101_001: DATA = 1'b0;
            15'b10111010_1101_010: DATA = 1'b0;
            15'b10111010_1101_011: DATA = 1'b0;
            15'b10111010_1101_100: DATA = 1'b0;
            15'b10111010_1101_101: DATA = 1'b0;
            15'b10111010_1101_110: DATA = 1'b0;
            15'b10111010_1101_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 3 Row 14
            15'b10111010_1110_000: DATA = 1'b0;
            15'b10111010_1110_001: DATA = 1'b0;
            15'b10111010_1110_010: DATA = 1'b0;
            15'b10111010_1110_011: DATA = 1'b0;
            15'b10111010_1110_100: DATA = 1'b0;
            15'b10111010_1110_101: DATA = 1'b0;
            15'b10111010_1110_110: DATA = 1'b0;
            15'b10111010_1110_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 3 Row 15
            15'b10111010_1111_000: DATA = 1'b0;
            15'b10111010_1111_001: DATA = 1'b0;
            15'b10111010_1111_010: DATA = 1'b0;
            15'b10111010_1111_011: DATA = 1'b0;
            15'b10111010_1111_100: DATA = 1'b0;
            15'b10111010_1111_101: DATA = 1'b0;
            15'b10111010_1111_110: DATA = 1'b0;
            15'b10111010_1111_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 4 Row 0
            15'b10111011_0000_000: DATA = 1'b0;
            15'b10111011_0000_001: DATA = 1'b0;
            15'b10111011_0000_010: DATA = 1'b0;
            15'b10111011_0000_011: DATA = 1'b0;
            15'b10111011_0000_100: DATA = 1'b0;
            15'b10111011_0000_101: DATA = 1'b0;
            15'b10111011_0000_110: DATA = 1'b0;
            15'b10111011_0000_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 4 Row 1
            15'b10111011_0001_000: DATA = 1'b0;
            15'b10111011_0001_001: DATA = 1'b0;
            15'b10111011_0001_010: DATA = 1'b0;
            15'b10111011_0001_011: DATA = 1'b0;
            15'b10111011_0001_100: DATA = 1'b0;
            15'b10111011_0001_101: DATA = 1'b0;
            15'b10111011_0001_110: DATA = 1'b0;
            15'b10111011_0001_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 4 Row 2
            15'b10111011_0010_000: DATA = 1'b0;
            15'b10111011_0010_001: DATA = 1'b0;
            15'b10111011_0010_010: DATA = 1'b0;
            15'b10111011_0010_011: DATA = 1'b0;
            15'b10111011_0010_100: DATA = 1'b0;
            15'b10111011_0010_101: DATA = 1'b0;
            15'b10111011_0010_110: DATA = 1'b0;
            15'b10111011_0010_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 4 Row 3
            15'b10111011_0011_000: DATA = 1'b0;
            15'b10111011_0011_001: DATA = 1'b0;
            15'b10111011_0011_010: DATA = 1'b0;
            15'b10111011_0011_011: DATA = 1'b0;
            15'b10111011_0011_100: DATA = 1'b0;
            15'b10111011_0011_101: DATA = 1'b0;
            15'b10111011_0011_110: DATA = 1'b0;
            15'b10111011_0011_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 4 Row 4
            15'b10111011_0100_000: DATA = 1'b0;
            15'b10111011_0100_001: DATA = 1'b0;
            15'b10111011_0100_010: DATA = 1'b0;
            15'b10111011_0100_011: DATA = 1'b0;
            15'b10111011_0100_100: DATA = 1'b0;
            15'b10111011_0100_101: DATA = 1'b0;
            15'b10111011_0100_110: DATA = 1'b0;
            15'b10111011_0100_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 4 Row 5
            15'b10111011_0101_000: DATA = 1'b0;
            15'b10111011_0101_001: DATA = 1'b0;
            15'b10111011_0101_010: DATA = 1'b0;
            15'b10111011_0101_011: DATA = 1'b0;
            15'b10111011_0101_100: DATA = 1'b0;
            15'b10111011_0101_101: DATA = 1'b0;
            15'b10111011_0101_110: DATA = 1'b0;
            15'b10111011_0101_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 4 Row 6
            15'b10111011_0110_000: DATA = 1'b0;
            15'b10111011_0110_001: DATA = 1'b0;
            15'b10111011_0110_010: DATA = 1'b0;
            15'b10111011_0110_011: DATA = 1'b0;
            15'b10111011_0110_100: DATA = 1'b0;
            15'b10111011_0110_101: DATA = 1'b0;
            15'b10111011_0110_110: DATA = 1'b0;
            15'b10111011_0110_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 4 Row 7
            15'b10111011_0111_000: DATA = 1'b0;
            15'b10111011_0111_001: DATA = 1'b0;
            15'b10111011_0111_010: DATA = 1'b0;
            15'b10111011_0111_011: DATA = 1'b0;
            15'b10111011_0111_100: DATA = 1'b0;
            15'b10111011_0111_101: DATA = 1'b0;
            15'b10111011_0111_110: DATA = 1'b0;
            15'b10111011_0111_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 4 Row 8
            15'b10111011_1000_000: DATA = 1'b0;
            15'b10111011_1000_001: DATA = 1'b0;
            15'b10111011_1000_010: DATA = 1'b0;
            15'b10111011_1000_011: DATA = 1'b0;
            15'b10111011_1000_100: DATA = 1'b0;
            15'b10111011_1000_101: DATA = 1'b0;
            15'b10111011_1000_110: DATA = 1'b0;
            15'b10111011_1000_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 4 Row 9
            15'b10111011_1001_000: DATA = 1'b0;
            15'b10111011_1001_001: DATA = 1'b0;
            15'b10111011_1001_010: DATA = 1'b0;
            15'b10111011_1001_011: DATA = 1'b0;
            15'b10111011_1001_100: DATA = 1'b0;
            15'b10111011_1001_101: DATA = 1'b0;
            15'b10111011_1001_110: DATA = 1'b0;
            15'b10111011_1001_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 4 Row 10
            15'b10111011_1010_000: DATA = 1'b0;
            15'b10111011_1010_001: DATA = 1'b0;
            15'b10111011_1010_010: DATA = 1'b0;
            15'b10111011_1010_011: DATA = 1'b0;
            15'b10111011_1010_100: DATA = 1'b0;
            15'b10111011_1010_101: DATA = 1'b0;
            15'b10111011_1010_110: DATA = 1'b0;
            15'b10111011_1010_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 4 Row 11
            15'b10111011_1011_000: DATA = 1'b0;
            15'b10111011_1011_001: DATA = 1'b0;
            15'b10111011_1011_010: DATA = 1'b0;
            15'b10111011_1011_011: DATA = 1'b0;
            15'b10111011_1011_100: DATA = 1'b0;
            15'b10111011_1011_101: DATA = 1'b0;
            15'b10111011_1011_110: DATA = 1'b0;
            15'b10111011_1011_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 4 Row 12
            15'b10111011_1100_000: DATA = 1'b0;
            15'b10111011_1100_001: DATA = 1'b0;
            15'b10111011_1100_010: DATA = 1'b0;
            15'b10111011_1100_011: DATA = 1'b0;
            15'b10111011_1100_100: DATA = 1'b0;
            15'b10111011_1100_101: DATA = 1'b0;
            15'b10111011_1100_110: DATA = 1'b0;
            15'b10111011_1100_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 4 Row 13
            15'b10111011_1101_000: DATA = 1'b0;
            15'b10111011_1101_001: DATA = 1'b0;
            15'b10111011_1101_010: DATA = 1'b0;
            15'b10111011_1101_011: DATA = 1'b0;
            15'b10111011_1101_100: DATA = 1'b0;
            15'b10111011_1101_101: DATA = 1'b0;
            15'b10111011_1101_110: DATA = 1'b0;
            15'b10111011_1101_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 4 Row 14
            15'b10111011_1110_000: DATA = 1'b0;
            15'b10111011_1110_001: DATA = 1'b0;
            15'b10111011_1110_010: DATA = 1'b0;
            15'b10111011_1110_011: DATA = 1'b0;
            15'b10111011_1110_100: DATA = 1'b0;
            15'b10111011_1110_101: DATA = 1'b0;
            15'b10111011_1110_110: DATA = 1'b0;
            15'b10111011_1110_111: DATA = 1'b0;
            // TRIANGLE- ROW 1 COL 4 Row 15
            15'b10111011_1111_000: DATA = 1'b0;
            15'b10111011_1111_001: DATA = 1'b0;
            15'b10111011_1111_010: DATA = 1'b0;
            15'b10111011_1111_011: DATA = 1'b0;
            15'b10111011_1111_100: DATA = 1'b0;
            15'b10111011_1111_101: DATA = 1'b0;
            15'b10111011_1111_110: DATA = 1'b0;
            15'b10111011_1111_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 0 Row 0
            15'b10111100_0000_000: DATA = 1'b0;
            15'b10111100_0000_001: DATA = 1'b0;
            15'b10111100_0000_010: DATA = 1'b0;
            15'b10111100_0000_011: DATA = 1'b0;
            15'b10111100_0000_100: DATA = 1'b0;
            15'b10111100_0000_101: DATA = 1'b0;
            15'b10111100_0000_110: DATA = 1'b0;
            15'b10111100_0000_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 0 Row 1
            15'b10111100_0001_000: DATA = 1'b0;
            15'b10111100_0001_001: DATA = 1'b0;
            15'b10111100_0001_010: DATA = 1'b0;
            15'b10111100_0001_011: DATA = 1'b0;
            15'b10111100_0001_100: DATA = 1'b0;
            15'b10111100_0001_101: DATA = 1'b0;
            15'b10111100_0001_110: DATA = 1'b0;
            15'b10111100_0001_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 0 Row 2
            15'b10111100_0010_000: DATA = 1'b0;
            15'b10111100_0010_001: DATA = 1'b0;
            15'b10111100_0010_010: DATA = 1'b0;
            15'b10111100_0010_011: DATA = 1'b0;
            15'b10111100_0010_100: DATA = 1'b0;
            15'b10111100_0010_101: DATA = 1'b0;
            15'b10111100_0010_110: DATA = 1'b0;
            15'b10111100_0010_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 0 Row 3
            15'b10111100_0011_000: DATA = 1'b0;
            15'b10111100_0011_001: DATA = 1'b0;
            15'b10111100_0011_010: DATA = 1'b0;
            15'b10111100_0011_011: DATA = 1'b0;
            15'b10111100_0011_100: DATA = 1'b0;
            15'b10111100_0011_101: DATA = 1'b0;
            15'b10111100_0011_110: DATA = 1'b0;
            15'b10111100_0011_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 0 Row 4
            15'b10111100_0100_000: DATA = 1'b0;
            15'b10111100_0100_001: DATA = 1'b0;
            15'b10111100_0100_010: DATA = 1'b0;
            15'b10111100_0100_011: DATA = 1'b0;
            15'b10111100_0100_100: DATA = 1'b0;
            15'b10111100_0100_101: DATA = 1'b0;
            15'b10111100_0100_110: DATA = 1'b0;
            15'b10111100_0100_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 0 Row 5
            15'b10111100_0101_000: DATA = 1'b0;
            15'b10111100_0101_001: DATA = 1'b0;
            15'b10111100_0101_010: DATA = 1'b0;
            15'b10111100_0101_011: DATA = 1'b0;
            15'b10111100_0101_100: DATA = 1'b0;
            15'b10111100_0101_101: DATA = 1'b0;
            15'b10111100_0101_110: DATA = 1'b0;
            15'b10111100_0101_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 0 Row 6
            15'b10111100_0110_000: DATA = 1'b0;
            15'b10111100_0110_001: DATA = 1'b0;
            15'b10111100_0110_010: DATA = 1'b0;
            15'b10111100_0110_011: DATA = 1'b0;
            15'b10111100_0110_100: DATA = 1'b0;
            15'b10111100_0110_101: DATA = 1'b0;
            15'b10111100_0110_110: DATA = 1'b0;
            15'b10111100_0110_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 0 Row 7
            15'b10111100_0111_000: DATA = 1'b0;
            15'b10111100_0111_001: DATA = 1'b0;
            15'b10111100_0111_010: DATA = 1'b0;
            15'b10111100_0111_011: DATA = 1'b0;
            15'b10111100_0111_100: DATA = 1'b0;
            15'b10111100_0111_101: DATA = 1'b0;
            15'b10111100_0111_110: DATA = 1'b0;
            15'b10111100_0111_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 0 Row 8
            15'b10111100_1000_000: DATA = 1'b0;
            15'b10111100_1000_001: DATA = 1'b0;
            15'b10111100_1000_010: DATA = 1'b0;
            15'b10111100_1000_011: DATA = 1'b0;
            15'b10111100_1000_100: DATA = 1'b0;
            15'b10111100_1000_101: DATA = 1'b0;
            15'b10111100_1000_110: DATA = 1'b0;
            15'b10111100_1000_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 0 Row 9
            15'b10111100_1001_000: DATA = 1'b0;
            15'b10111100_1001_001: DATA = 1'b0;
            15'b10111100_1001_010: DATA = 1'b0;
            15'b10111100_1001_011: DATA = 1'b0;
            15'b10111100_1001_100: DATA = 1'b0;
            15'b10111100_1001_101: DATA = 1'b0;
            15'b10111100_1001_110: DATA = 1'b0;
            15'b10111100_1001_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 0 Row 10
            15'b10111100_1010_000: DATA = 1'b0;
            15'b10111100_1010_001: DATA = 1'b0;
            15'b10111100_1010_010: DATA = 1'b0;
            15'b10111100_1010_011: DATA = 1'b0;
            15'b10111100_1010_100: DATA = 1'b0;
            15'b10111100_1010_101: DATA = 1'b0;
            15'b10111100_1010_110: DATA = 1'b0;
            15'b10111100_1010_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 0 Row 11
            15'b10111100_1011_000: DATA = 1'b0;
            15'b10111100_1011_001: DATA = 1'b0;
            15'b10111100_1011_010: DATA = 1'b0;
            15'b10111100_1011_011: DATA = 1'b0;
            15'b10111100_1011_100: DATA = 1'b0;
            15'b10111100_1011_101: DATA = 1'b0;
            15'b10111100_1011_110: DATA = 1'b0;
            15'b10111100_1011_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 0 Row 12
            15'b10111100_1100_000: DATA = 1'b0;
            15'b10111100_1100_001: DATA = 1'b0;
            15'b10111100_1100_010: DATA = 1'b0;
            15'b10111100_1100_011: DATA = 1'b0;
            15'b10111100_1100_100: DATA = 1'b0;
            15'b10111100_1100_101: DATA = 1'b0;
            15'b10111100_1100_110: DATA = 1'b0;
            15'b10111100_1100_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 0 Row 13
            15'b10111100_1101_000: DATA = 1'b0;
            15'b10111100_1101_001: DATA = 1'b0;
            15'b10111100_1101_010: DATA = 1'b0;
            15'b10111100_1101_011: DATA = 1'b0;
            15'b10111100_1101_100: DATA = 1'b0;
            15'b10111100_1101_101: DATA = 1'b0;
            15'b10111100_1101_110: DATA = 1'b0;
            15'b10111100_1101_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 0 Row 14
            15'b10111100_1110_000: DATA = 1'b0;
            15'b10111100_1110_001: DATA = 1'b0;
            15'b10111100_1110_010: DATA = 1'b0;
            15'b10111100_1110_011: DATA = 1'b0;
            15'b10111100_1110_100: DATA = 1'b0;
            15'b10111100_1110_101: DATA = 1'b0;
            15'b10111100_1110_110: DATA = 1'b0;
            15'b10111100_1110_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 0 Row 15
            15'b10111100_1111_000: DATA = 1'b0;
            15'b10111100_1111_001: DATA = 1'b0;
            15'b10111100_1111_010: DATA = 1'b0;
            15'b10111100_1111_011: DATA = 1'b0;
            15'b10111100_1111_100: DATA = 1'b0;
            15'b10111100_1111_101: DATA = 1'b0;
            15'b10111100_1111_110: DATA = 1'b0;
            15'b10111100_1111_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 1 Row 0
            15'b10111101_0000_000: DATA = 1'b0;
            15'b10111101_0000_001: DATA = 1'b0;
            15'b10111101_0000_010: DATA = 1'b0;
            15'b10111101_0000_011: DATA = 1'b0;
            15'b10111101_0000_100: DATA = 1'b0;
            15'b10111101_0000_101: DATA = 1'b0;
            15'b10111101_0000_110: DATA = 1'b0;
            15'b10111101_0000_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 1 Row 1
            15'b10111101_0001_000: DATA = 1'b0;
            15'b10111101_0001_001: DATA = 1'b0;
            15'b10111101_0001_010: DATA = 1'b0;
            15'b10111101_0001_011: DATA = 1'b0;
            15'b10111101_0001_100: DATA = 1'b0;
            15'b10111101_0001_101: DATA = 1'b0;
            15'b10111101_0001_110: DATA = 1'b0;
            15'b10111101_0001_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 1 Row 2
            15'b10111101_0010_000: DATA = 1'b0;
            15'b10111101_0010_001: DATA = 1'b0;
            15'b10111101_0010_010: DATA = 1'b0;
            15'b10111101_0010_011: DATA = 1'b0;
            15'b10111101_0010_100: DATA = 1'b0;
            15'b10111101_0010_101: DATA = 1'b0;
            15'b10111101_0010_110: DATA = 1'b0;
            15'b10111101_0010_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 1 Row 3
            15'b10111101_0011_000: DATA = 1'b0;
            15'b10111101_0011_001: DATA = 1'b0;
            15'b10111101_0011_010: DATA = 1'b0;
            15'b10111101_0011_011: DATA = 1'b0;
            15'b10111101_0011_100: DATA = 1'b0;
            15'b10111101_0011_101: DATA = 1'b0;
            15'b10111101_0011_110: DATA = 1'b0;
            15'b10111101_0011_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 1 Row 4
            15'b10111101_0100_000: DATA = 1'b0;
            15'b10111101_0100_001: DATA = 1'b0;
            15'b10111101_0100_010: DATA = 1'b0;
            15'b10111101_0100_011: DATA = 1'b0;
            15'b10111101_0100_100: DATA = 1'b0;
            15'b10111101_0100_101: DATA = 1'b0;
            15'b10111101_0100_110: DATA = 1'b0;
            15'b10111101_0100_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 1 Row 5
            15'b10111101_0101_000: DATA = 1'b0;
            15'b10111101_0101_001: DATA = 1'b0;
            15'b10111101_0101_010: DATA = 1'b0;
            15'b10111101_0101_011: DATA = 1'b0;
            15'b10111101_0101_100: DATA = 1'b0;
            15'b10111101_0101_101: DATA = 1'b0;
            15'b10111101_0101_110: DATA = 1'b0;
            15'b10111101_0101_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 1 Row 6
            15'b10111101_0110_000: DATA = 1'b0;
            15'b10111101_0110_001: DATA = 1'b0;
            15'b10111101_0110_010: DATA = 1'b0;
            15'b10111101_0110_011: DATA = 1'b0;
            15'b10111101_0110_100: DATA = 1'b0;
            15'b10111101_0110_101: DATA = 1'b0;
            15'b10111101_0110_110: DATA = 1'b0;
            15'b10111101_0110_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 1 Row 7
            15'b10111101_0111_000: DATA = 1'b0;
            15'b10111101_0111_001: DATA = 1'b0;
            15'b10111101_0111_010: DATA = 1'b0;
            15'b10111101_0111_011: DATA = 1'b0;
            15'b10111101_0111_100: DATA = 1'b0;
            15'b10111101_0111_101: DATA = 1'b0;
            15'b10111101_0111_110: DATA = 1'b0;
            15'b10111101_0111_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 1 Row 8
            15'b10111101_1000_000: DATA = 1'b0;
            15'b10111101_1000_001: DATA = 1'b0;
            15'b10111101_1000_010: DATA = 1'b0;
            15'b10111101_1000_011: DATA = 1'b0;
            15'b10111101_1000_100: DATA = 1'b0;
            15'b10111101_1000_101: DATA = 1'b0;
            15'b10111101_1000_110: DATA = 1'b0;
            15'b10111101_1000_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 1 Row 9
            15'b10111101_1001_000: DATA = 1'b0;
            15'b10111101_1001_001: DATA = 1'b0;
            15'b10111101_1001_010: DATA = 1'b0;
            15'b10111101_1001_011: DATA = 1'b0;
            15'b10111101_1001_100: DATA = 1'b0;
            15'b10111101_1001_101: DATA = 1'b0;
            15'b10111101_1001_110: DATA = 1'b0;
            15'b10111101_1001_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 1 Row 10
            15'b10111101_1010_000: DATA = 1'b0;
            15'b10111101_1010_001: DATA = 1'b0;
            15'b10111101_1010_010: DATA = 1'b0;
            15'b10111101_1010_011: DATA = 1'b0;
            15'b10111101_1010_100: DATA = 1'b0;
            15'b10111101_1010_101: DATA = 1'b0;
            15'b10111101_1010_110: DATA = 1'b0;
            15'b10111101_1010_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 1 Row 11
            15'b10111101_1011_000: DATA = 1'b0;
            15'b10111101_1011_001: DATA = 1'b0;
            15'b10111101_1011_010: DATA = 1'b0;
            15'b10111101_1011_011: DATA = 1'b0;
            15'b10111101_1011_100: DATA = 1'b0;
            15'b10111101_1011_101: DATA = 1'b0;
            15'b10111101_1011_110: DATA = 1'b0;
            15'b10111101_1011_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 1 Row 12
            15'b10111101_1100_000: DATA = 1'b0;
            15'b10111101_1100_001: DATA = 1'b0;
            15'b10111101_1100_010: DATA = 1'b0;
            15'b10111101_1100_011: DATA = 1'b0;
            15'b10111101_1100_100: DATA = 1'b0;
            15'b10111101_1100_101: DATA = 1'b0;
            15'b10111101_1100_110: DATA = 1'b0;
            15'b10111101_1100_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 1 Row 13
            15'b10111101_1101_000: DATA = 1'b0;
            15'b10111101_1101_001: DATA = 1'b0;
            15'b10111101_1101_010: DATA = 1'b0;
            15'b10111101_1101_011: DATA = 1'b0;
            15'b10111101_1101_100: DATA = 1'b0;
            15'b10111101_1101_101: DATA = 1'b0;
            15'b10111101_1101_110: DATA = 1'b0;
            15'b10111101_1101_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 1 Row 14
            15'b10111101_1110_000: DATA = 1'b0;
            15'b10111101_1110_001: DATA = 1'b0;
            15'b10111101_1110_010: DATA = 1'b0;
            15'b10111101_1110_011: DATA = 1'b0;
            15'b10111101_1110_100: DATA = 1'b0;
            15'b10111101_1110_101: DATA = 1'b0;
            15'b10111101_1110_110: DATA = 1'b0;
            15'b10111101_1110_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 1 Row 15
            15'b10111101_1111_000: DATA = 1'b0;
            15'b10111101_1111_001: DATA = 1'b0;
            15'b10111101_1111_010: DATA = 1'b0;
            15'b10111101_1111_011: DATA = 1'b0;
            15'b10111101_1111_100: DATA = 1'b0;
            15'b10111101_1111_101: DATA = 1'b0;
            15'b10111101_1111_110: DATA = 1'b0;
            15'b10111101_1111_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 2 Row 0
            15'b10111110_0000_000: DATA = 1'b0;
            15'b10111110_0000_001: DATA = 1'b0;
            15'b10111110_0000_010: DATA = 1'b0;
            15'b10111110_0000_011: DATA = 1'b0;
            15'b10111110_0000_100: DATA = 1'b0;
            15'b10111110_0000_101: DATA = 1'b0;
            15'b10111110_0000_110: DATA = 1'b0;
            15'b10111110_0000_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 2 Row 1
            15'b10111110_0001_000: DATA = 1'b0;
            15'b10111110_0001_001: DATA = 1'b0;
            15'b10111110_0001_010: DATA = 1'b0;
            15'b10111110_0001_011: DATA = 1'b0;
            15'b10111110_0001_100: DATA = 1'b0;
            15'b10111110_0001_101: DATA = 1'b0;
            15'b10111110_0001_110: DATA = 1'b0;
            15'b10111110_0001_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 2 Row 2
            15'b10111110_0010_000: DATA = 1'b0;
            15'b10111110_0010_001: DATA = 1'b0;
            15'b10111110_0010_010: DATA = 1'b0;
            15'b10111110_0010_011: DATA = 1'b0;
            15'b10111110_0010_100: DATA = 1'b0;
            15'b10111110_0010_101: DATA = 1'b0;
            15'b10111110_0010_110: DATA = 1'b0;
            15'b10111110_0010_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 2 Row 3
            15'b10111110_0011_000: DATA = 1'b0;
            15'b10111110_0011_001: DATA = 1'b0;
            15'b10111110_0011_010: DATA = 1'b0;
            15'b10111110_0011_011: DATA = 1'b0;
            15'b10111110_0011_100: DATA = 1'b0;
            15'b10111110_0011_101: DATA = 1'b0;
            15'b10111110_0011_110: DATA = 1'b0;
            15'b10111110_0011_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 2 Row 4
            15'b10111110_0100_000: DATA = 1'b0;
            15'b10111110_0100_001: DATA = 1'b0;
            15'b10111110_0100_010: DATA = 1'b0;
            15'b10111110_0100_011: DATA = 1'b0;
            15'b10111110_0100_100: DATA = 1'b0;
            15'b10111110_0100_101: DATA = 1'b0;
            15'b10111110_0100_110: DATA = 1'b0;
            15'b10111110_0100_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 2 Row 5
            15'b10111110_0101_000: DATA = 1'b0;
            15'b10111110_0101_001: DATA = 1'b0;
            15'b10111110_0101_010: DATA = 1'b0;
            15'b10111110_0101_011: DATA = 1'b0;
            15'b10111110_0101_100: DATA = 1'b0;
            15'b10111110_0101_101: DATA = 1'b0;
            15'b10111110_0101_110: DATA = 1'b0;
            15'b10111110_0101_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 2 Row 6
            15'b10111110_0110_000: DATA = 1'b0;
            15'b10111110_0110_001: DATA = 1'b0;
            15'b10111110_0110_010: DATA = 1'b0;
            15'b10111110_0110_011: DATA = 1'b0;
            15'b10111110_0110_100: DATA = 1'b0;
            15'b10111110_0110_101: DATA = 1'b0;
            15'b10111110_0110_110: DATA = 1'b0;
            15'b10111110_0110_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 2 Row 7
            15'b10111110_0111_000: DATA = 1'b0;
            15'b10111110_0111_001: DATA = 1'b0;
            15'b10111110_0111_010: DATA = 1'b0;
            15'b10111110_0111_011: DATA = 1'b0;
            15'b10111110_0111_100: DATA = 1'b0;
            15'b10111110_0111_101: DATA = 1'b0;
            15'b10111110_0111_110: DATA = 1'b0;
            15'b10111110_0111_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 2 Row 8
            15'b10111110_1000_000: DATA = 1'b0;
            15'b10111110_1000_001: DATA = 1'b0;
            15'b10111110_1000_010: DATA = 1'b0;
            15'b10111110_1000_011: DATA = 1'b0;
            15'b10111110_1000_100: DATA = 1'b0;
            15'b10111110_1000_101: DATA = 1'b0;
            15'b10111110_1000_110: DATA = 1'b0;
            15'b10111110_1000_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 2 Row 9
            15'b10111110_1001_000: DATA = 1'b0;
            15'b10111110_1001_001: DATA = 1'b0;
            15'b10111110_1001_010: DATA = 1'b0;
            15'b10111110_1001_011: DATA = 1'b0;
            15'b10111110_1001_100: DATA = 1'b0;
            15'b10111110_1001_101: DATA = 1'b0;
            15'b10111110_1001_110: DATA = 1'b0;
            15'b10111110_1001_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 2 Row 10
            15'b10111110_1010_000: DATA = 1'b0;
            15'b10111110_1010_001: DATA = 1'b0;
            15'b10111110_1010_010: DATA = 1'b0;
            15'b10111110_1010_011: DATA = 1'b0;
            15'b10111110_1010_100: DATA = 1'b0;
            15'b10111110_1010_101: DATA = 1'b0;
            15'b10111110_1010_110: DATA = 1'b0;
            15'b10111110_1010_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 2 Row 11
            15'b10111110_1011_000: DATA = 1'b0;
            15'b10111110_1011_001: DATA = 1'b0;
            15'b10111110_1011_010: DATA = 1'b0;
            15'b10111110_1011_011: DATA = 1'b0;
            15'b10111110_1011_100: DATA = 1'b0;
            15'b10111110_1011_101: DATA = 1'b0;
            15'b10111110_1011_110: DATA = 1'b0;
            15'b10111110_1011_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 0 COL 2 Row 12
            15'b10111110_1100_000: DATA = 1'b0;
            15'b10111110_1100_001: DATA = 1'b0;
            15'b10111110_1100_010: DATA = 1'b0;
            15'b10111110_1100_011: DATA = 1'b0;
            15'b10111110_1100_100: DATA = 1'b0;
            15'b10111110_1100_101: DATA = 1'b0;
            15'b10111110_1100_110: DATA = 1'b1;
            15'b10111110_1100_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 0 COL 2 Row 13
            15'b10111110_1101_000: DATA = 1'b0;
            15'b10111110_1101_001: DATA = 1'b0;
            15'b10111110_1101_010: DATA = 1'b0;
            15'b10111110_1101_011: DATA = 1'b0;
            15'b10111110_1101_100: DATA = 1'b0;
            15'b10111110_1101_101: DATA = 1'b1;
            15'b10111110_1101_110: DATA = 1'b1;
            15'b10111110_1101_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 2 Row 14
            15'b10111110_1110_000: DATA = 1'b0;
            15'b10111110_1110_001: DATA = 1'b0;
            15'b10111110_1110_010: DATA = 1'b0;
            15'b10111110_1110_011: DATA = 1'b0;
            15'b10111110_1110_100: DATA = 1'b1;
            15'b10111110_1110_101: DATA = 1'b1;
            15'b10111110_1110_110: DATA = 1'b0;
            15'b10111110_1110_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 2 Row 15
            15'b10111110_1111_000: DATA = 1'b0;
            15'b10111110_1111_001: DATA = 1'b0;
            15'b10111110_1111_010: DATA = 1'b1;
            15'b10111110_1111_011: DATA = 1'b1;
            15'b10111110_1111_100: DATA = 1'b1;
            15'b10111110_1111_101: DATA = 1'b0;
            15'b10111110_1111_110: DATA = 1'b0;
            15'b10111110_1111_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 3 Row 0
            15'b10111111_0000_000: DATA = 1'b0;
            15'b10111111_0000_001: DATA = 1'b0;
            15'b10111111_0000_010: DATA = 1'b0;
            15'b10111111_0000_011: DATA = 1'b0;
            15'b10111111_0000_100: DATA = 1'b0;
            15'b10111111_0000_101: DATA = 1'b0;
            15'b10111111_0000_110: DATA = 1'b0;
            15'b10111111_0000_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 3 Row 1
            15'b10111111_0001_000: DATA = 1'b0;
            15'b10111111_0001_001: DATA = 1'b0;
            15'b10111111_0001_010: DATA = 1'b0;
            15'b10111111_0001_011: DATA = 1'b0;
            15'b10111111_0001_100: DATA = 1'b0;
            15'b10111111_0001_101: DATA = 1'b0;
            15'b10111111_0001_110: DATA = 1'b0;
            15'b10111111_0001_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 3 Row 2
            15'b10111111_0010_000: DATA = 1'b0;
            15'b10111111_0010_001: DATA = 1'b0;
            15'b10111111_0010_010: DATA = 1'b0;
            15'b10111111_0010_011: DATA = 1'b0;
            15'b10111111_0010_100: DATA = 1'b0;
            15'b10111111_0010_101: DATA = 1'b0;
            15'b10111111_0010_110: DATA = 1'b0;
            15'b10111111_0010_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 3 Row 3
            15'b10111111_0011_000: DATA = 1'b0;
            15'b10111111_0011_001: DATA = 1'b0;
            15'b10111111_0011_010: DATA = 1'b0;
            15'b10111111_0011_011: DATA = 1'b0;
            15'b10111111_0011_100: DATA = 1'b0;
            15'b10111111_0011_101: DATA = 1'b0;
            15'b10111111_0011_110: DATA = 1'b0;
            15'b10111111_0011_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 3 Row 4
            15'b10111111_0100_000: DATA = 1'b0;
            15'b10111111_0100_001: DATA = 1'b0;
            15'b10111111_0100_010: DATA = 1'b0;
            15'b10111111_0100_011: DATA = 1'b0;
            15'b10111111_0100_100: DATA = 1'b0;
            15'b10111111_0100_101: DATA = 1'b0;
            15'b10111111_0100_110: DATA = 1'b0;
            15'b10111111_0100_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 3 Row 5
            15'b10111111_0101_000: DATA = 1'b0;
            15'b10111111_0101_001: DATA = 1'b0;
            15'b10111111_0101_010: DATA = 1'b0;
            15'b10111111_0101_011: DATA = 1'b0;
            15'b10111111_0101_100: DATA = 1'b0;
            15'b10111111_0101_101: DATA = 1'b0;
            15'b10111111_0101_110: DATA = 1'b0;
            15'b10111111_0101_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 0 COL 3 Row 6
            15'b10111111_0110_000: DATA = 1'b0;
            15'b10111111_0110_001: DATA = 1'b0;
            15'b10111111_0110_010: DATA = 1'b0;
            15'b10111111_0110_011: DATA = 1'b0;
            15'b10111111_0110_100: DATA = 1'b0;
            15'b10111111_0110_101: DATA = 1'b0;
            15'b10111111_0110_110: DATA = 1'b1;
            15'b10111111_0110_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 0 COL 3 Row 7
            15'b10111111_0111_000: DATA = 1'b0;
            15'b10111111_0111_001: DATA = 1'b0;
            15'b10111111_0111_010: DATA = 1'b0;
            15'b10111111_0111_011: DATA = 1'b0;
            15'b10111111_0111_100: DATA = 1'b1;
            15'b10111111_0111_101: DATA = 1'b1;
            15'b10111111_0111_110: DATA = 1'b1;
            15'b10111111_0111_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 3 Row 8
            15'b10111111_1000_000: DATA = 1'b0;
            15'b10111111_1000_001: DATA = 1'b0;
            15'b10111111_1000_010: DATA = 1'b0;
            15'b10111111_1000_011: DATA = 1'b1;
            15'b10111111_1000_100: DATA = 1'b1;
            15'b10111111_1000_101: DATA = 1'b0;
            15'b10111111_1000_110: DATA = 1'b0;
            15'b10111111_1000_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 3 Row 9
            15'b10111111_1001_000: DATA = 1'b0;
            15'b10111111_1001_001: DATA = 1'b0;
            15'b10111111_1001_010: DATA = 1'b1;
            15'b10111111_1001_011: DATA = 1'b1;
            15'b10111111_1001_100: DATA = 1'b0;
            15'b10111111_1001_101: DATA = 1'b0;
            15'b10111111_1001_110: DATA = 1'b0;
            15'b10111111_1001_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 3 Row 10
            15'b10111111_1010_000: DATA = 1'b0;
            15'b10111111_1010_001: DATA = 1'b1;
            15'b10111111_1010_010: DATA = 1'b1;
            15'b10111111_1010_011: DATA = 1'b0;
            15'b10111111_1010_100: DATA = 1'b0;
            15'b10111111_1010_101: DATA = 1'b0;
            15'b10111111_1010_110: DATA = 1'b0;
            15'b10111111_1010_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 3 Row 11
            15'b10111111_1011_000: DATA = 1'b1;
            15'b10111111_1011_001: DATA = 1'b1;
            15'b10111111_1011_010: DATA = 1'b0;
            15'b10111111_1011_011: DATA = 1'b0;
            15'b10111111_1011_100: DATA = 1'b0;
            15'b10111111_1011_101: DATA = 1'b0;
            15'b10111111_1011_110: DATA = 1'b0;
            15'b10111111_1011_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 3 Row 12
            15'b10111111_1100_000: DATA = 1'b0;
            15'b10111111_1100_001: DATA = 1'b0;
            15'b10111111_1100_010: DATA = 1'b0;
            15'b10111111_1100_011: DATA = 1'b0;
            15'b10111111_1100_100: DATA = 1'b0;
            15'b10111111_1100_101: DATA = 1'b0;
            15'b10111111_1100_110: DATA = 1'b0;
            15'b10111111_1100_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 3 Row 13
            15'b10111111_1101_000: DATA = 1'b0;
            15'b10111111_1101_001: DATA = 1'b0;
            15'b10111111_1101_010: DATA = 1'b0;
            15'b10111111_1101_011: DATA = 1'b0;
            15'b10111111_1101_100: DATA = 1'b0;
            15'b10111111_1101_101: DATA = 1'b0;
            15'b10111111_1101_110: DATA = 1'b0;
            15'b10111111_1101_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 3 Row 14
            15'b10111111_1110_000: DATA = 1'b0;
            15'b10111111_1110_001: DATA = 1'b0;
            15'b10111111_1110_010: DATA = 1'b0;
            15'b10111111_1110_011: DATA = 1'b0;
            15'b10111111_1110_100: DATA = 1'b0;
            15'b10111111_1110_101: DATA = 1'b0;
            15'b10111111_1110_110: DATA = 1'b0;
            15'b10111111_1110_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 3 Row 15
            15'b10111111_1111_000: DATA = 1'b0;
            15'b10111111_1111_001: DATA = 1'b0;
            15'b10111111_1111_010: DATA = 1'b0;
            15'b10111111_1111_011: DATA = 1'b0;
            15'b10111111_1111_100: DATA = 1'b0;
            15'b10111111_1111_101: DATA = 1'b0;
            15'b10111111_1111_110: DATA = 1'b0;
            15'b10111111_1111_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 0 COL 4 Row 0
            15'b11000000_0000_000: DATA = 1'b0;
            15'b11000000_0000_001: DATA = 1'b0;
            15'b11000000_0000_010: DATA = 1'b0;
            15'b11000000_0000_011: DATA = 1'b0;
            15'b11000000_0000_100: DATA = 1'b0;
            15'b11000000_0000_101: DATA = 1'b0;
            15'b11000000_0000_110: DATA = 1'b1;
            15'b11000000_0000_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 0 COL 4 Row 1
            15'b11000000_0001_000: DATA = 1'b0;
            15'b11000000_0001_001: DATA = 1'b0;
            15'b11000000_0001_010: DATA = 1'b0;
            15'b11000000_0001_011: DATA = 1'b0;
            15'b11000000_0001_100: DATA = 1'b1;
            15'b11000000_0001_101: DATA = 1'b1;
            15'b11000000_0001_110: DATA = 1'b0;
            15'b11000000_0001_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 0 COL 4 Row 2
            15'b11000000_0010_000: DATA = 1'b0;
            15'b11000000_0010_001: DATA = 1'b0;
            15'b11000000_0010_010: DATA = 1'b0;
            15'b11000000_0010_011: DATA = 1'b1;
            15'b11000000_0010_100: DATA = 1'b1;
            15'b11000000_0010_101: DATA = 1'b0;
            15'b11000000_0010_110: DATA = 1'b0;
            15'b11000000_0010_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 0 COL 4 Row 3
            15'b11000000_0011_000: DATA = 1'b0;
            15'b11000000_0011_001: DATA = 1'b1;
            15'b11000000_0011_010: DATA = 1'b1;
            15'b11000000_0011_011: DATA = 1'b1;
            15'b11000000_0011_100: DATA = 1'b0;
            15'b11000000_0011_101: DATA = 1'b0;
            15'b11000000_0011_110: DATA = 1'b0;
            15'b11000000_0011_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 0 COL 4 Row 4
            15'b11000000_0100_000: DATA = 1'b1;
            15'b11000000_0100_001: DATA = 1'b1;
            15'b11000000_0100_010: DATA = 1'b0;
            15'b11000000_0100_011: DATA = 1'b0;
            15'b11000000_0100_100: DATA = 1'b0;
            15'b11000000_0100_101: DATA = 1'b0;
            15'b11000000_0100_110: DATA = 1'b0;
            15'b11000000_0100_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 0 COL 4 Row 5
            15'b11000000_0101_000: DATA = 1'b1;
            15'b11000000_0101_001: DATA = 1'b0;
            15'b11000000_0101_010: DATA = 1'b0;
            15'b11000000_0101_011: DATA = 1'b0;
            15'b11000000_0101_100: DATA = 1'b0;
            15'b11000000_0101_101: DATA = 1'b0;
            15'b11000000_0101_110: DATA = 1'b0;
            15'b11000000_0101_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 0 COL 4 Row 6
            15'b11000000_0110_000: DATA = 1'b0;
            15'b11000000_0110_001: DATA = 1'b0;
            15'b11000000_0110_010: DATA = 1'b0;
            15'b11000000_0110_011: DATA = 1'b0;
            15'b11000000_0110_100: DATA = 1'b0;
            15'b11000000_0110_101: DATA = 1'b0;
            15'b11000000_0110_110: DATA = 1'b0;
            15'b11000000_0110_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 0 COL 4 Row 7
            15'b11000000_0111_000: DATA = 1'b0;
            15'b11000000_0111_001: DATA = 1'b0;
            15'b11000000_0111_010: DATA = 1'b0;
            15'b11000000_0111_011: DATA = 1'b0;
            15'b11000000_0111_100: DATA = 1'b0;
            15'b11000000_0111_101: DATA = 1'b0;
            15'b11000000_0111_110: DATA = 1'b0;
            15'b11000000_0111_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 0 COL 4 Row 8
            15'b11000000_1000_000: DATA = 1'b0;
            15'b11000000_1000_001: DATA = 1'b0;
            15'b11000000_1000_010: DATA = 1'b0;
            15'b11000000_1000_011: DATA = 1'b0;
            15'b11000000_1000_100: DATA = 1'b0;
            15'b11000000_1000_101: DATA = 1'b0;
            15'b11000000_1000_110: DATA = 1'b0;
            15'b11000000_1000_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 0 COL 4 Row 9
            15'b11000000_1001_000: DATA = 1'b0;
            15'b11000000_1001_001: DATA = 1'b0;
            15'b11000000_1001_010: DATA = 1'b0;
            15'b11000000_1001_011: DATA = 1'b0;
            15'b11000000_1001_100: DATA = 1'b0;
            15'b11000000_1001_101: DATA = 1'b0;
            15'b11000000_1001_110: DATA = 1'b0;
            15'b11000000_1001_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 0 COL 4 Row 10
            15'b11000000_1010_000: DATA = 1'b0;
            15'b11000000_1010_001: DATA = 1'b0;
            15'b11000000_1010_010: DATA = 1'b0;
            15'b11000000_1010_011: DATA = 1'b0;
            15'b11000000_1010_100: DATA = 1'b0;
            15'b11000000_1010_101: DATA = 1'b0;
            15'b11000000_1010_110: DATA = 1'b0;
            15'b11000000_1010_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 0 COL 4 Row 11
            15'b11000000_1011_000: DATA = 1'b0;
            15'b11000000_1011_001: DATA = 1'b0;
            15'b11000000_1011_010: DATA = 1'b0;
            15'b11000000_1011_011: DATA = 1'b0;
            15'b11000000_1011_100: DATA = 1'b0;
            15'b11000000_1011_101: DATA = 1'b0;
            15'b11000000_1011_110: DATA = 1'b0;
            15'b11000000_1011_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 0 COL 4 Row 12
            15'b11000000_1100_000: DATA = 1'b0;
            15'b11000000_1100_001: DATA = 1'b0;
            15'b11000000_1100_010: DATA = 1'b0;
            15'b11000000_1100_011: DATA = 1'b0;
            15'b11000000_1100_100: DATA = 1'b0;
            15'b11000000_1100_101: DATA = 1'b0;
            15'b11000000_1100_110: DATA = 1'b0;
            15'b11000000_1100_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 0 COL 4 Row 13
            15'b11000000_1101_000: DATA = 1'b0;
            15'b11000000_1101_001: DATA = 1'b0;
            15'b11000000_1101_010: DATA = 1'b0;
            15'b11000000_1101_011: DATA = 1'b0;
            15'b11000000_1101_100: DATA = 1'b0;
            15'b11000000_1101_101: DATA = 1'b0;
            15'b11000000_1101_110: DATA = 1'b0;
            15'b11000000_1101_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 0 COL 4 Row 14
            15'b11000000_1110_000: DATA = 1'b0;
            15'b11000000_1110_001: DATA = 1'b0;
            15'b11000000_1110_010: DATA = 1'b0;
            15'b11000000_1110_011: DATA = 1'b0;
            15'b11000000_1110_100: DATA = 1'b0;
            15'b11000000_1110_101: DATA = 1'b0;
            15'b11000000_1110_110: DATA = 1'b0;
            15'b11000000_1110_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 0 COL 4 Row 15
            15'b11000000_1111_000: DATA = 1'b0;
            15'b11000000_1111_001: DATA = 1'b0;
            15'b11000000_1111_010: DATA = 1'b0;
            15'b11000000_1111_011: DATA = 1'b0;
            15'b11000000_1111_100: DATA = 1'b0;
            15'b11000000_1111_101: DATA = 1'b0;
            15'b11000000_1111_110: DATA = 1'b0;
            15'b11000000_1111_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 1 COL 0 Row 0
            15'b11000001_0000_000: DATA = 1'b0;
            15'b11000001_0000_001: DATA = 1'b0;
            15'b11000001_0000_010: DATA = 1'b0;
            15'b11000001_0000_011: DATA = 1'b0;
            15'b11000001_0000_100: DATA = 1'b0;
            15'b11000001_0000_101: DATA = 1'b0;
            15'b11000001_0000_110: DATA = 1'b0;
            15'b11000001_0000_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 0 Row 1
            15'b11000001_0001_000: DATA = 1'b0;
            15'b11000001_0001_001: DATA = 1'b0;
            15'b11000001_0001_010: DATA = 1'b0;
            15'b11000001_0001_011: DATA = 1'b0;
            15'b11000001_0001_100: DATA = 1'b0;
            15'b11000001_0001_101: DATA = 1'b0;
            15'b11000001_0001_110: DATA = 1'b0;
            15'b11000001_0001_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 0 Row 2
            15'b11000001_0010_000: DATA = 1'b0;
            15'b11000001_0010_001: DATA = 1'b0;
            15'b11000001_0010_010: DATA = 1'b0;
            15'b11000001_0010_011: DATA = 1'b0;
            15'b11000001_0010_100: DATA = 1'b0;
            15'b11000001_0010_101: DATA = 1'b0;
            15'b11000001_0010_110: DATA = 1'b0;
            15'b11000001_0010_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 0 Row 3
            15'b11000001_0011_000: DATA = 1'b0;
            15'b11000001_0011_001: DATA = 1'b0;
            15'b11000001_0011_010: DATA = 1'b0;
            15'b11000001_0011_011: DATA = 1'b0;
            15'b11000001_0011_100: DATA = 1'b0;
            15'b11000001_0011_101: DATA = 1'b0;
            15'b11000001_0011_110: DATA = 1'b0;
            15'b11000001_0011_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 0 Row 4
            15'b11000001_0100_000: DATA = 1'b0;
            15'b11000001_0100_001: DATA = 1'b0;
            15'b11000001_0100_010: DATA = 1'b0;
            15'b11000001_0100_011: DATA = 1'b0;
            15'b11000001_0100_100: DATA = 1'b0;
            15'b11000001_0100_101: DATA = 1'b0;
            15'b11000001_0100_110: DATA = 1'b0;
            15'b11000001_0100_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 0 Row 5
            15'b11000001_0101_000: DATA = 1'b0;
            15'b11000001_0101_001: DATA = 1'b0;
            15'b11000001_0101_010: DATA = 1'b0;
            15'b11000001_0101_011: DATA = 1'b0;
            15'b11000001_0101_100: DATA = 1'b0;
            15'b11000001_0101_101: DATA = 1'b0;
            15'b11000001_0101_110: DATA = 1'b0;
            15'b11000001_0101_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 0 Row 6
            15'b11000001_0110_000: DATA = 1'b0;
            15'b11000001_0110_001: DATA = 1'b0;
            15'b11000001_0110_010: DATA = 1'b0;
            15'b11000001_0110_011: DATA = 1'b0;
            15'b11000001_0110_100: DATA = 1'b0;
            15'b11000001_0110_101: DATA = 1'b0;
            15'b11000001_0110_110: DATA = 1'b0;
            15'b11000001_0110_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 0 Row 7
            15'b11000001_0111_000: DATA = 1'b0;
            15'b11000001_0111_001: DATA = 1'b0;
            15'b11000001_0111_010: DATA = 1'b0;
            15'b11000001_0111_011: DATA = 1'b0;
            15'b11000001_0111_100: DATA = 1'b0;
            15'b11000001_0111_101: DATA = 1'b0;
            15'b11000001_0111_110: DATA = 1'b0;
            15'b11000001_0111_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 0 Row 8
            15'b11000001_1000_000: DATA = 1'b0;
            15'b11000001_1000_001: DATA = 1'b0;
            15'b11000001_1000_010: DATA = 1'b0;
            15'b11000001_1000_011: DATA = 1'b0;
            15'b11000001_1000_100: DATA = 1'b0;
            15'b11000001_1000_101: DATA = 1'b0;
            15'b11000001_1000_110: DATA = 1'b0;
            15'b11000001_1000_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 1 COL 0 Row 9
            15'b11000001_1001_000: DATA = 1'b0;
            15'b11000001_1001_001: DATA = 1'b0;
            15'b11000001_1001_010: DATA = 1'b0;
            15'b11000001_1001_011: DATA = 1'b0;
            15'b11000001_1001_100: DATA = 1'b0;
            15'b11000001_1001_101: DATA = 1'b0;
            15'b11000001_1001_110: DATA = 1'b1;
            15'b11000001_1001_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 1 COL 0 Row 10
            15'b11000001_1010_000: DATA = 1'b0;
            15'b11000001_1010_001: DATA = 1'b0;
            15'b11000001_1010_010: DATA = 1'b0;
            15'b11000001_1010_011: DATA = 1'b0;
            15'b11000001_1010_100: DATA = 1'b0;
            15'b11000001_1010_101: DATA = 1'b1;
            15'b11000001_1010_110: DATA = 1'b1;
            15'b11000001_1010_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 0 Row 11
            15'b11000001_1011_000: DATA = 1'b0;
            15'b11000001_1011_001: DATA = 1'b0;
            15'b11000001_1011_010: DATA = 1'b0;
            15'b11000001_1011_011: DATA = 1'b1;
            15'b11000001_1011_100: DATA = 1'b1;
            15'b11000001_1011_101: DATA = 1'b1;
            15'b11000001_1011_110: DATA = 1'b0;
            15'b11000001_1011_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 0 Row 12
            15'b11000001_1100_000: DATA = 1'b0;
            15'b11000001_1100_001: DATA = 1'b0;
            15'b11000001_1100_010: DATA = 1'b1;
            15'b11000001_1100_011: DATA = 1'b1;
            15'b11000001_1100_100: DATA = 1'b0;
            15'b11000001_1100_101: DATA = 1'b0;
            15'b11000001_1100_110: DATA = 1'b0;
            15'b11000001_1100_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 0 Row 13
            15'b11000001_1101_000: DATA = 1'b0;
            15'b11000001_1101_001: DATA = 1'b1;
            15'b11000001_1101_010: DATA = 1'b1;
            15'b11000001_1101_011: DATA = 1'b0;
            15'b11000001_1101_100: DATA = 1'b0;
            15'b11000001_1101_101: DATA = 1'b0;
            15'b11000001_1101_110: DATA = 1'b0;
            15'b11000001_1101_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 0 Row 14
            15'b11000001_1110_000: DATA = 1'b1;
            15'b11000001_1110_001: DATA = 1'b1;
            15'b11000001_1110_010: DATA = 1'b0;
            15'b11000001_1110_011: DATA = 1'b0;
            15'b11000001_1110_100: DATA = 1'b0;
            15'b11000001_1110_101: DATA = 1'b0;
            15'b11000001_1110_110: DATA = 1'b0;
            15'b11000001_1110_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 0 Row 15
            15'b11000001_1111_000: DATA = 1'b1;
            15'b11000001_1111_001: DATA = 1'b0;
            15'b11000001_1111_010: DATA = 1'b0;
            15'b11000001_1111_011: DATA = 1'b0;
            15'b11000001_1111_100: DATA = 1'b0;
            15'b11000001_1111_101: DATA = 1'b0;
            15'b11000001_1111_110: DATA = 1'b0;
            15'b11000001_1111_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 1 Row 0
            15'b11000010_0000_000: DATA = 1'b0;
            15'b11000010_0000_001: DATA = 1'b0;
            15'b11000010_0000_010: DATA = 1'b0;
            15'b11000010_0000_011: DATA = 1'b0;
            15'b11000010_0000_100: DATA = 1'b0;
            15'b11000010_0000_101: DATA = 1'b0;
            15'b11000010_0000_110: DATA = 1'b0;
            15'b11000010_0000_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 1 Row 1
            15'b11000010_0001_000: DATA = 1'b0;
            15'b11000010_0001_001: DATA = 1'b0;
            15'b11000010_0001_010: DATA = 1'b0;
            15'b11000010_0001_011: DATA = 1'b0;
            15'b11000010_0001_100: DATA = 1'b0;
            15'b11000010_0001_101: DATA = 1'b0;
            15'b11000010_0001_110: DATA = 1'b0;
            15'b11000010_0001_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 1 Row 2
            15'b11000010_0010_000: DATA = 1'b0;
            15'b11000010_0010_001: DATA = 1'b0;
            15'b11000010_0010_010: DATA = 1'b0;
            15'b11000010_0010_011: DATA = 1'b0;
            15'b11000010_0010_100: DATA = 1'b0;
            15'b11000010_0010_101: DATA = 1'b0;
            15'b11000010_0010_110: DATA = 1'b0;
            15'b11000010_0010_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 1 COL 1 Row 3
            15'b11000010_0011_000: DATA = 1'b0;
            15'b11000010_0011_001: DATA = 1'b0;
            15'b11000010_0011_010: DATA = 1'b0;
            15'b11000010_0011_011: DATA = 1'b0;
            15'b11000010_0011_100: DATA = 1'b0;
            15'b11000010_0011_101: DATA = 1'b1;
            15'b11000010_0011_110: DATA = 1'b1;
            15'b11000010_0011_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 1 COL 1 Row 4
            15'b11000010_0100_000: DATA = 1'b0;
            15'b11000010_0100_001: DATA = 1'b0;
            15'b11000010_0100_010: DATA = 1'b0;
            15'b11000010_0100_011: DATA = 1'b0;
            15'b11000010_0100_100: DATA = 1'b1;
            15'b11000010_0100_101: DATA = 1'b1;
            15'b11000010_0100_110: DATA = 1'b0;
            15'b11000010_0100_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 1 Row 5
            15'b11000010_0101_000: DATA = 1'b0;
            15'b11000010_0101_001: DATA = 1'b0;
            15'b11000010_0101_010: DATA = 1'b0;
            15'b11000010_0101_011: DATA = 1'b1;
            15'b11000010_0101_100: DATA = 1'b1;
            15'b11000010_0101_101: DATA = 1'b0;
            15'b11000010_0101_110: DATA = 1'b0;
            15'b11000010_0101_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 1 Row 6
            15'b11000010_0110_000: DATA = 1'b0;
            15'b11000010_0110_001: DATA = 1'b0;
            15'b11000010_0110_010: DATA = 1'b1;
            15'b11000010_0110_011: DATA = 1'b1;
            15'b11000010_0110_100: DATA = 1'b0;
            15'b11000010_0110_101: DATA = 1'b0;
            15'b11000010_0110_110: DATA = 1'b0;
            15'b11000010_0110_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 1 Row 7
            15'b11000010_0111_000: DATA = 1'b1;
            15'b11000010_0111_001: DATA = 1'b1;
            15'b11000010_0111_010: DATA = 1'b1;
            15'b11000010_0111_011: DATA = 1'b0;
            15'b11000010_0111_100: DATA = 1'b0;
            15'b11000010_0111_101: DATA = 1'b0;
            15'b11000010_0111_110: DATA = 1'b0;
            15'b11000010_0111_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 1 Row 8
            15'b11000010_1000_000: DATA = 1'b1;
            15'b11000010_1000_001: DATA = 1'b0;
            15'b11000010_1000_010: DATA = 1'b0;
            15'b11000010_1000_011: DATA = 1'b0;
            15'b11000010_1000_100: DATA = 1'b0;
            15'b11000010_1000_101: DATA = 1'b0;
            15'b11000010_1000_110: DATA = 1'b0;
            15'b11000010_1000_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 1 Row 9
            15'b11000010_1001_000: DATA = 1'b0;
            15'b11000010_1001_001: DATA = 1'b0;
            15'b11000010_1001_010: DATA = 1'b0;
            15'b11000010_1001_011: DATA = 1'b0;
            15'b11000010_1001_100: DATA = 1'b0;
            15'b11000010_1001_101: DATA = 1'b0;
            15'b11000010_1001_110: DATA = 1'b0;
            15'b11000010_1001_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 1 Row 10
            15'b11000010_1010_000: DATA = 1'b0;
            15'b11000010_1010_001: DATA = 1'b0;
            15'b11000010_1010_010: DATA = 1'b0;
            15'b11000010_1010_011: DATA = 1'b0;
            15'b11000010_1010_100: DATA = 1'b0;
            15'b11000010_1010_101: DATA = 1'b0;
            15'b11000010_1010_110: DATA = 1'b0;
            15'b11000010_1010_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 1 Row 11
            15'b11000010_1011_000: DATA = 1'b0;
            15'b11000010_1011_001: DATA = 1'b0;
            15'b11000010_1011_010: DATA = 1'b0;
            15'b11000010_1011_011: DATA = 1'b0;
            15'b11000010_1011_100: DATA = 1'b0;
            15'b11000010_1011_101: DATA = 1'b0;
            15'b11000010_1011_110: DATA = 1'b0;
            15'b11000010_1011_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 1 Row 12
            15'b11000010_1100_000: DATA = 1'b0;
            15'b11000010_1100_001: DATA = 1'b0;
            15'b11000010_1100_010: DATA = 1'b0;
            15'b11000010_1100_011: DATA = 1'b0;
            15'b11000010_1100_100: DATA = 1'b0;
            15'b11000010_1100_101: DATA = 1'b0;
            15'b11000010_1100_110: DATA = 1'b0;
            15'b11000010_1100_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 1 Row 13
            15'b11000010_1101_000: DATA = 1'b0;
            15'b11000010_1101_001: DATA = 1'b0;
            15'b11000010_1101_010: DATA = 1'b0;
            15'b11000010_1101_011: DATA = 1'b0;
            15'b11000010_1101_100: DATA = 1'b0;
            15'b11000010_1101_101: DATA = 1'b0;
            15'b11000010_1101_110: DATA = 1'b0;
            15'b11000010_1101_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 1 Row 14
            15'b11000010_1110_000: DATA = 1'b0;
            15'b11000010_1110_001: DATA = 1'b0;
            15'b11000010_1110_010: DATA = 1'b0;
            15'b11000010_1110_011: DATA = 1'b0;
            15'b11000010_1110_100: DATA = 1'b0;
            15'b11000010_1110_101: DATA = 1'b0;
            15'b11000010_1110_110: DATA = 1'b0;
            15'b11000010_1110_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 1 Row 15
            15'b11000010_1111_000: DATA = 1'b0;
            15'b11000010_1111_001: DATA = 1'b0;
            15'b11000010_1111_010: DATA = 1'b0;
            15'b11000010_1111_011: DATA = 1'b0;
            15'b11000010_1111_100: DATA = 1'b0;
            15'b11000010_1111_101: DATA = 1'b0;
            15'b11000010_1111_110: DATA = 1'b0;
            15'b11000010_1111_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 2 Row 0
            15'b11000011_0000_000: DATA = 1'b0;
            15'b11000011_0000_001: DATA = 1'b1;
            15'b11000011_0000_010: DATA = 1'b1;
            15'b11000011_0000_011: DATA = 1'b0;
            15'b11000011_0000_100: DATA = 1'b0;
            15'b11000011_0000_101: DATA = 1'b0;
            15'b11000011_0000_110: DATA = 1'b0;
            15'b11000011_0000_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 2 Row 1
            15'b11000011_0001_000: DATA = 1'b1;
            15'b11000011_0001_001: DATA = 1'b1;
            15'b11000011_0001_010: DATA = 1'b0;
            15'b11000011_0001_011: DATA = 1'b0;
            15'b11000011_0001_100: DATA = 1'b0;
            15'b11000011_0001_101: DATA = 1'b0;
            15'b11000011_0001_110: DATA = 1'b0;
            15'b11000011_0001_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 2 Row 2
            15'b11000011_0010_000: DATA = 1'b1;
            15'b11000011_0010_001: DATA = 1'b0;
            15'b11000011_0010_010: DATA = 1'b0;
            15'b11000011_0010_011: DATA = 1'b0;
            15'b11000011_0010_100: DATA = 1'b0;
            15'b11000011_0010_101: DATA = 1'b0;
            15'b11000011_0010_110: DATA = 1'b0;
            15'b11000011_0010_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 2 Row 3
            15'b11000011_0011_000: DATA = 1'b0;
            15'b11000011_0011_001: DATA = 1'b0;
            15'b11000011_0011_010: DATA = 1'b0;
            15'b11000011_0011_011: DATA = 1'b0;
            15'b11000011_0011_100: DATA = 1'b0;
            15'b11000011_0011_101: DATA = 1'b0;
            15'b11000011_0011_110: DATA = 1'b0;
            15'b11000011_0011_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 2 Row 4
            15'b11000011_0100_000: DATA = 1'b0;
            15'b11000011_0100_001: DATA = 1'b0;
            15'b11000011_0100_010: DATA = 1'b0;
            15'b11000011_0100_011: DATA = 1'b0;
            15'b11000011_0100_100: DATA = 1'b0;
            15'b11000011_0100_101: DATA = 1'b0;
            15'b11000011_0100_110: DATA = 1'b0;
            15'b11000011_0100_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 2 Row 5
            15'b11000011_0101_000: DATA = 1'b0;
            15'b11000011_0101_001: DATA = 1'b0;
            15'b11000011_0101_010: DATA = 1'b0;
            15'b11000011_0101_011: DATA = 1'b0;
            15'b11000011_0101_100: DATA = 1'b0;
            15'b11000011_0101_101: DATA = 1'b0;
            15'b11000011_0101_110: DATA = 1'b0;
            15'b11000011_0101_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 2 Row 6
            15'b11000011_0110_000: DATA = 1'b0;
            15'b11000011_0110_001: DATA = 1'b0;
            15'b11000011_0110_010: DATA = 1'b0;
            15'b11000011_0110_011: DATA = 1'b0;
            15'b11000011_0110_100: DATA = 1'b0;
            15'b11000011_0110_101: DATA = 1'b0;
            15'b11000011_0110_110: DATA = 1'b0;
            15'b11000011_0110_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 2 Row 7
            15'b11000011_0111_000: DATA = 1'b0;
            15'b11000011_0111_001: DATA = 1'b0;
            15'b11000011_0111_010: DATA = 1'b0;
            15'b11000011_0111_011: DATA = 1'b0;
            15'b11000011_0111_100: DATA = 1'b0;
            15'b11000011_0111_101: DATA = 1'b0;
            15'b11000011_0111_110: DATA = 1'b0;
            15'b11000011_0111_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 2 Row 8
            15'b11000011_1000_000: DATA = 1'b0;
            15'b11000011_1000_001: DATA = 1'b0;
            15'b11000011_1000_010: DATA = 1'b0;
            15'b11000011_1000_011: DATA = 1'b0;
            15'b11000011_1000_100: DATA = 1'b0;
            15'b11000011_1000_101: DATA = 1'b0;
            15'b11000011_1000_110: DATA = 1'b0;
            15'b11000011_1000_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 2 Row 9
            15'b11000011_1001_000: DATA = 1'b0;
            15'b11000011_1001_001: DATA = 1'b0;
            15'b11000011_1001_010: DATA = 1'b0;
            15'b11000011_1001_011: DATA = 1'b0;
            15'b11000011_1001_100: DATA = 1'b0;
            15'b11000011_1001_101: DATA = 1'b0;
            15'b11000011_1001_110: DATA = 1'b0;
            15'b11000011_1001_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 2 Row 10
            15'b11000011_1010_000: DATA = 1'b0;
            15'b11000011_1010_001: DATA = 1'b0;
            15'b11000011_1010_010: DATA = 1'b0;
            15'b11000011_1010_011: DATA = 1'b0;
            15'b11000011_1010_100: DATA = 1'b0;
            15'b11000011_1010_101: DATA = 1'b0;
            15'b11000011_1010_110: DATA = 1'b0;
            15'b11000011_1010_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 2 Row 11
            15'b11000011_1011_000: DATA = 1'b0;
            15'b11000011_1011_001: DATA = 1'b0;
            15'b11000011_1011_010: DATA = 1'b0;
            15'b11000011_1011_011: DATA = 1'b0;
            15'b11000011_1011_100: DATA = 1'b0;
            15'b11000011_1011_101: DATA = 1'b0;
            15'b11000011_1011_110: DATA = 1'b0;
            15'b11000011_1011_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 2 Row 12
            15'b11000011_1100_000: DATA = 1'b0;
            15'b11000011_1100_001: DATA = 1'b0;
            15'b11000011_1100_010: DATA = 1'b0;
            15'b11000011_1100_011: DATA = 1'b0;
            15'b11000011_1100_100: DATA = 1'b0;
            15'b11000011_1100_101: DATA = 1'b0;
            15'b11000011_1100_110: DATA = 1'b0;
            15'b11000011_1100_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 2 Row 13
            15'b11000011_1101_000: DATA = 1'b0;
            15'b11000011_1101_001: DATA = 1'b0;
            15'b11000011_1101_010: DATA = 1'b0;
            15'b11000011_1101_011: DATA = 1'b0;
            15'b11000011_1101_100: DATA = 1'b0;
            15'b11000011_1101_101: DATA = 1'b0;
            15'b11000011_1101_110: DATA = 1'b0;
            15'b11000011_1101_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 2 Row 14
            15'b11000011_1110_000: DATA = 1'b0;
            15'b11000011_1110_001: DATA = 1'b0;
            15'b11000011_1110_010: DATA = 1'b0;
            15'b11000011_1110_011: DATA = 1'b0;
            15'b11000011_1110_100: DATA = 1'b0;
            15'b11000011_1110_101: DATA = 1'b0;
            15'b11000011_1110_110: DATA = 1'b0;
            15'b11000011_1110_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 2 Row 15
            15'b11000011_1111_000: DATA = 1'b0;
            15'b11000011_1111_001: DATA = 1'b0;
            15'b11000011_1111_010: DATA = 1'b0;
            15'b11000011_1111_011: DATA = 1'b0;
            15'b11000011_1111_100: DATA = 1'b0;
            15'b11000011_1111_101: DATA = 1'b0;
            15'b11000011_1111_110: DATA = 1'b0;
            15'b11000011_1111_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 3 Row 0
            15'b11000100_0000_000: DATA = 1'b0;
            15'b11000100_0000_001: DATA = 1'b0;
            15'b11000100_0000_010: DATA = 1'b0;
            15'b11000100_0000_011: DATA = 1'b0;
            15'b11000100_0000_100: DATA = 1'b0;
            15'b11000100_0000_101: DATA = 1'b0;
            15'b11000100_0000_110: DATA = 1'b0;
            15'b11000100_0000_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 3 Row 1
            15'b11000100_0001_000: DATA = 1'b0;
            15'b11000100_0001_001: DATA = 1'b0;
            15'b11000100_0001_010: DATA = 1'b0;
            15'b11000100_0001_011: DATA = 1'b0;
            15'b11000100_0001_100: DATA = 1'b0;
            15'b11000100_0001_101: DATA = 1'b0;
            15'b11000100_0001_110: DATA = 1'b0;
            15'b11000100_0001_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 3 Row 2
            15'b11000100_0010_000: DATA = 1'b0;
            15'b11000100_0010_001: DATA = 1'b0;
            15'b11000100_0010_010: DATA = 1'b0;
            15'b11000100_0010_011: DATA = 1'b0;
            15'b11000100_0010_100: DATA = 1'b0;
            15'b11000100_0010_101: DATA = 1'b0;
            15'b11000100_0010_110: DATA = 1'b0;
            15'b11000100_0010_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 3 Row 3
            15'b11000100_0011_000: DATA = 1'b0;
            15'b11000100_0011_001: DATA = 1'b0;
            15'b11000100_0011_010: DATA = 1'b0;
            15'b11000100_0011_011: DATA = 1'b0;
            15'b11000100_0011_100: DATA = 1'b0;
            15'b11000100_0011_101: DATA = 1'b0;
            15'b11000100_0011_110: DATA = 1'b0;
            15'b11000100_0011_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 3 Row 4
            15'b11000100_0100_000: DATA = 1'b0;
            15'b11000100_0100_001: DATA = 1'b0;
            15'b11000100_0100_010: DATA = 1'b0;
            15'b11000100_0100_011: DATA = 1'b0;
            15'b11000100_0100_100: DATA = 1'b0;
            15'b11000100_0100_101: DATA = 1'b0;
            15'b11000100_0100_110: DATA = 1'b0;
            15'b11000100_0100_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 3 Row 5
            15'b11000100_0101_000: DATA = 1'b0;
            15'b11000100_0101_001: DATA = 1'b0;
            15'b11000100_0101_010: DATA = 1'b0;
            15'b11000100_0101_011: DATA = 1'b0;
            15'b11000100_0101_100: DATA = 1'b0;
            15'b11000100_0101_101: DATA = 1'b0;
            15'b11000100_0101_110: DATA = 1'b0;
            15'b11000100_0101_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 3 Row 6
            15'b11000100_0110_000: DATA = 1'b0;
            15'b11000100_0110_001: DATA = 1'b0;
            15'b11000100_0110_010: DATA = 1'b0;
            15'b11000100_0110_011: DATA = 1'b0;
            15'b11000100_0110_100: DATA = 1'b0;
            15'b11000100_0110_101: DATA = 1'b0;
            15'b11000100_0110_110: DATA = 1'b0;
            15'b11000100_0110_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 3 Row 7
            15'b11000100_0111_000: DATA = 1'b0;
            15'b11000100_0111_001: DATA = 1'b0;
            15'b11000100_0111_010: DATA = 1'b0;
            15'b11000100_0111_011: DATA = 1'b0;
            15'b11000100_0111_100: DATA = 1'b0;
            15'b11000100_0111_101: DATA = 1'b0;
            15'b11000100_0111_110: DATA = 1'b0;
            15'b11000100_0111_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 3 Row 8
            15'b11000100_1000_000: DATA = 1'b0;
            15'b11000100_1000_001: DATA = 1'b0;
            15'b11000100_1000_010: DATA = 1'b0;
            15'b11000100_1000_011: DATA = 1'b0;
            15'b11000100_1000_100: DATA = 1'b0;
            15'b11000100_1000_101: DATA = 1'b0;
            15'b11000100_1000_110: DATA = 1'b0;
            15'b11000100_1000_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 3 Row 9
            15'b11000100_1001_000: DATA = 1'b0;
            15'b11000100_1001_001: DATA = 1'b0;
            15'b11000100_1001_010: DATA = 1'b0;
            15'b11000100_1001_011: DATA = 1'b0;
            15'b11000100_1001_100: DATA = 1'b0;
            15'b11000100_1001_101: DATA = 1'b0;
            15'b11000100_1001_110: DATA = 1'b0;
            15'b11000100_1001_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 3 Row 10
            15'b11000100_1010_000: DATA = 1'b0;
            15'b11000100_1010_001: DATA = 1'b0;
            15'b11000100_1010_010: DATA = 1'b0;
            15'b11000100_1010_011: DATA = 1'b0;
            15'b11000100_1010_100: DATA = 1'b0;
            15'b11000100_1010_101: DATA = 1'b0;
            15'b11000100_1010_110: DATA = 1'b0;
            15'b11000100_1010_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 3 Row 11
            15'b11000100_1011_000: DATA = 1'b0;
            15'b11000100_1011_001: DATA = 1'b0;
            15'b11000100_1011_010: DATA = 1'b0;
            15'b11000100_1011_011: DATA = 1'b0;
            15'b11000100_1011_100: DATA = 1'b0;
            15'b11000100_1011_101: DATA = 1'b0;
            15'b11000100_1011_110: DATA = 1'b0;
            15'b11000100_1011_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 3 Row 12
            15'b11000100_1100_000: DATA = 1'b0;
            15'b11000100_1100_001: DATA = 1'b0;
            15'b11000100_1100_010: DATA = 1'b0;
            15'b11000100_1100_011: DATA = 1'b0;
            15'b11000100_1100_100: DATA = 1'b0;
            15'b11000100_1100_101: DATA = 1'b0;
            15'b11000100_1100_110: DATA = 1'b0;
            15'b11000100_1100_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 3 Row 13
            15'b11000100_1101_000: DATA = 1'b0;
            15'b11000100_1101_001: DATA = 1'b0;
            15'b11000100_1101_010: DATA = 1'b0;
            15'b11000100_1101_011: DATA = 1'b0;
            15'b11000100_1101_100: DATA = 1'b0;
            15'b11000100_1101_101: DATA = 1'b0;
            15'b11000100_1101_110: DATA = 1'b0;
            15'b11000100_1101_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 3 Row 14
            15'b11000100_1110_000: DATA = 1'b0;
            15'b11000100_1110_001: DATA = 1'b0;
            15'b11000100_1110_010: DATA = 1'b0;
            15'b11000100_1110_011: DATA = 1'b0;
            15'b11000100_1110_100: DATA = 1'b0;
            15'b11000100_1110_101: DATA = 1'b0;
            15'b11000100_1110_110: DATA = 1'b0;
            15'b11000100_1110_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 3 Row 15
            15'b11000100_1111_000: DATA = 1'b0;
            15'b11000100_1111_001: DATA = 1'b0;
            15'b11000100_1111_010: DATA = 1'b0;
            15'b11000100_1111_011: DATA = 1'b0;
            15'b11000100_1111_100: DATA = 1'b0;
            15'b11000100_1111_101: DATA = 1'b0;
            15'b11000100_1111_110: DATA = 1'b0;
            15'b11000100_1111_111: DATA = 1'b0;
            //SAWTOOTH+ ROW 1 COL 4 Row 0
            15'b11000101_0000_000: DATA = 1'b0;
            15'b11000101_0000_001: DATA = 1'b0;
            15'b11000101_0000_010: DATA = 1'b0;
            15'b11000101_0000_011: DATA = 1'b0;
            15'b11000101_0000_100: DATA = 1'b0;
            15'b11000101_0000_101: DATA = 1'b0;
            15'b11000101_0000_110: DATA = 1'b0;
            15'b11000101_0000_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 1 COL 4 Row 1
            15'b11000101_0001_000: DATA = 1'b0;
            15'b11000101_0001_001: DATA = 1'b0;
            15'b11000101_0001_010: DATA = 1'b0;
            15'b11000101_0001_011: DATA = 1'b0;
            15'b11000101_0001_100: DATA = 1'b0;
            15'b11000101_0001_101: DATA = 1'b0;
            15'b11000101_0001_110: DATA = 1'b0;
            15'b11000101_0001_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 1 COL 4 Row 2
            15'b11000101_0010_000: DATA = 1'b0;
            15'b11000101_0010_001: DATA = 1'b0;
            15'b11000101_0010_010: DATA = 1'b0;
            15'b11000101_0010_011: DATA = 1'b0;
            15'b11000101_0010_100: DATA = 1'b0;
            15'b11000101_0010_101: DATA = 1'b0;
            15'b11000101_0010_110: DATA = 1'b0;
            15'b11000101_0010_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 1 COL 4 Row 3
            15'b11000101_0011_000: DATA = 1'b0;
            15'b11000101_0011_001: DATA = 1'b0;
            15'b11000101_0011_010: DATA = 1'b0;
            15'b11000101_0011_011: DATA = 1'b0;
            15'b11000101_0011_100: DATA = 1'b0;
            15'b11000101_0011_101: DATA = 1'b0;
            15'b11000101_0011_110: DATA = 1'b0;
            15'b11000101_0011_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 1 COL 4 Row 4
            15'b11000101_0100_000: DATA = 1'b0;
            15'b11000101_0100_001: DATA = 1'b0;
            15'b11000101_0100_010: DATA = 1'b0;
            15'b11000101_0100_011: DATA = 1'b0;
            15'b11000101_0100_100: DATA = 1'b0;
            15'b11000101_0100_101: DATA = 1'b0;
            15'b11000101_0100_110: DATA = 1'b0;
            15'b11000101_0100_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 1 COL 4 Row 5
            15'b11000101_0101_000: DATA = 1'b0;
            15'b11000101_0101_001: DATA = 1'b0;
            15'b11000101_0101_010: DATA = 1'b0;
            15'b11000101_0101_011: DATA = 1'b0;
            15'b11000101_0101_100: DATA = 1'b0;
            15'b11000101_0101_101: DATA = 1'b0;
            15'b11000101_0101_110: DATA = 1'b0;
            15'b11000101_0101_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 1 COL 4 Row 6
            15'b11000101_0110_000: DATA = 1'b0;
            15'b11000101_0110_001: DATA = 1'b0;
            15'b11000101_0110_010: DATA = 1'b0;
            15'b11000101_0110_011: DATA = 1'b0;
            15'b11000101_0110_100: DATA = 1'b0;
            15'b11000101_0110_101: DATA = 1'b0;
            15'b11000101_0110_110: DATA = 1'b0;
            15'b11000101_0110_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 1 COL 4 Row 7
            15'b11000101_0111_000: DATA = 1'b0;
            15'b11000101_0111_001: DATA = 1'b0;
            15'b11000101_0111_010: DATA = 1'b0;
            15'b11000101_0111_011: DATA = 1'b0;
            15'b11000101_0111_100: DATA = 1'b0;
            15'b11000101_0111_101: DATA = 1'b0;
            15'b11000101_0111_110: DATA = 1'b0;
            15'b11000101_0111_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 1 COL 4 Row 8
            15'b11000101_1000_000: DATA = 1'b0;
            15'b11000101_1000_001: DATA = 1'b0;
            15'b11000101_1000_010: DATA = 1'b0;
            15'b11000101_1000_011: DATA = 1'b0;
            15'b11000101_1000_100: DATA = 1'b0;
            15'b11000101_1000_101: DATA = 1'b0;
            15'b11000101_1000_110: DATA = 1'b0;
            15'b11000101_1000_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 1 COL 4 Row 9
            15'b11000101_1001_000: DATA = 1'b0;
            15'b11000101_1001_001: DATA = 1'b0;
            15'b11000101_1001_010: DATA = 1'b0;
            15'b11000101_1001_011: DATA = 1'b0;
            15'b11000101_1001_100: DATA = 1'b0;
            15'b11000101_1001_101: DATA = 1'b0;
            15'b11000101_1001_110: DATA = 1'b0;
            15'b11000101_1001_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 1 COL 4 Row 10
            15'b11000101_1010_000: DATA = 1'b0;
            15'b11000101_1010_001: DATA = 1'b0;
            15'b11000101_1010_010: DATA = 1'b0;
            15'b11000101_1010_011: DATA = 1'b0;
            15'b11000101_1010_100: DATA = 1'b0;
            15'b11000101_1010_101: DATA = 1'b0;
            15'b11000101_1010_110: DATA = 1'b0;
            15'b11000101_1010_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 1 COL 4 Row 11
            15'b11000101_1011_000: DATA = 1'b0;
            15'b11000101_1011_001: DATA = 1'b0;
            15'b11000101_1011_010: DATA = 1'b0;
            15'b11000101_1011_011: DATA = 1'b0;
            15'b11000101_1011_100: DATA = 1'b0;
            15'b11000101_1011_101: DATA = 1'b0;
            15'b11000101_1011_110: DATA = 1'b0;
            15'b11000101_1011_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 1 COL 4 Row 12
            15'b11000101_1100_000: DATA = 1'b0;
            15'b11000101_1100_001: DATA = 1'b0;
            15'b11000101_1100_010: DATA = 1'b0;
            15'b11000101_1100_011: DATA = 1'b0;
            15'b11000101_1100_100: DATA = 1'b0;
            15'b11000101_1100_101: DATA = 1'b0;
            15'b11000101_1100_110: DATA = 1'b0;
            15'b11000101_1100_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 1 COL 4 Row 13
            15'b11000101_1101_000: DATA = 1'b0;
            15'b11000101_1101_001: DATA = 1'b0;
            15'b11000101_1101_010: DATA = 1'b0;
            15'b11000101_1101_011: DATA = 1'b0;
            15'b11000101_1101_100: DATA = 1'b0;
            15'b11000101_1101_101: DATA = 1'b0;
            15'b11000101_1101_110: DATA = 1'b0;
            15'b11000101_1101_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 1 COL 4 Row 14
            15'b11000101_1110_000: DATA = 1'b0;
            15'b11000101_1110_001: DATA = 1'b0;
            15'b11000101_1110_010: DATA = 1'b0;
            15'b11000101_1110_011: DATA = 1'b0;
            15'b11000101_1110_100: DATA = 1'b0;
            15'b11000101_1110_101: DATA = 1'b0;
            15'b11000101_1110_110: DATA = 1'b0;
            15'b11000101_1110_111: DATA = 1'b1;
            //SAWTOOTH+ ROW 1 COL 4 Row 15
            15'b11000101_1111_000: DATA = 1'b0;
            15'b11000101_1111_001: DATA = 1'b0;
            15'b11000101_1111_010: DATA = 1'b0;
            15'b11000101_1111_011: DATA = 1'b0;
            15'b11000101_1111_100: DATA = 1'b0;
            15'b11000101_1111_101: DATA = 1'b0;
            15'b11000101_1111_110: DATA = 1'b0;
            15'b11000101_1111_111: DATA = 1'b1;
            //VERTICAL LEFT 0 COL 0 Row 0
            15'b11000110_0000_000: DATA = 1'b1;
            15'b11000110_0000_001: DATA = 1'b0;
            15'b11000110_0000_010: DATA = 1'b0;
            15'b11000110_0000_011: DATA = 1'b0;
            15'b11000110_0000_100: DATA = 1'b0;
            15'b11000110_0000_101: DATA = 1'b0;
            15'b11000110_0000_110: DATA = 1'b0;
            15'b11000110_0000_111: DATA = 1'b0;
            //VERTICAL LEFT 0 COL 0 Row 1
            15'b11000110_0001_000: DATA = 1'b1;
            15'b11000110_0001_001: DATA = 1'b0;
            15'b11000110_0001_010: DATA = 1'b0;
            15'b11000110_0001_011: DATA = 1'b0;
            15'b11000110_0001_100: DATA = 1'b0;
            15'b11000110_0001_101: DATA = 1'b0;
            15'b11000110_0001_110: DATA = 1'b0;
            15'b11000110_0001_111: DATA = 1'b0;
            //VERTICAL LEFT 0 COL 0 Row 2
            15'b11000110_0010_000: DATA = 1'b1;
            15'b11000110_0010_001: DATA = 1'b0;
            15'b11000110_0010_010: DATA = 1'b0;
            15'b11000110_0010_011: DATA = 1'b0;
            15'b11000110_0010_100: DATA = 1'b0;
            15'b11000110_0010_101: DATA = 1'b0;
            15'b11000110_0010_110: DATA = 1'b0;
            15'b11000110_0010_111: DATA = 1'b0;
            //VERTICAL LEFT 0 COL 0 Row 3
            15'b11000110_0011_000: DATA = 1'b1;
            15'b11000110_0011_001: DATA = 1'b0;
            15'b11000110_0011_010: DATA = 1'b0;
            15'b11000110_0011_011: DATA = 1'b0;
            15'b11000110_0011_100: DATA = 1'b0;
            15'b11000110_0011_101: DATA = 1'b0;
            15'b11000110_0011_110: DATA = 1'b0;
            15'b11000110_0011_111: DATA = 1'b0;
            //VERTICAL LEFT 0 COL 0 Row 4
            15'b11000110_0100_000: DATA = 1'b1;
            15'b11000110_0100_001: DATA = 1'b0;
            15'b11000110_0100_010: DATA = 1'b0;
            15'b11000110_0100_011: DATA = 1'b0;
            15'b11000110_0100_100: DATA = 1'b0;
            15'b11000110_0100_101: DATA = 1'b0;
            15'b11000110_0100_110: DATA = 1'b0;
            15'b11000110_0100_111: DATA = 1'b0;
            //VERTICAL LEFT 0 COL 0 Row 5
            15'b11000110_0101_000: DATA = 1'b1;
            15'b11000110_0101_001: DATA = 1'b0;
            15'b11000110_0101_010: DATA = 1'b0;
            15'b11000110_0101_011: DATA = 1'b0;
            15'b11000110_0101_100: DATA = 1'b0;
            15'b11000110_0101_101: DATA = 1'b0;
            15'b11000110_0101_110: DATA = 1'b0;
            15'b11000110_0101_111: DATA = 1'b0;
            //VERTICAL LEFT 0 COL 0 Row 6
            15'b11000110_0110_000: DATA = 1'b1;
            15'b11000110_0110_001: DATA = 1'b0;
            15'b11000110_0110_010: DATA = 1'b0;
            15'b11000110_0110_011: DATA = 1'b0;
            15'b11000110_0110_100: DATA = 1'b0;
            15'b11000110_0110_101: DATA = 1'b0;
            15'b11000110_0110_110: DATA = 1'b0;
            15'b11000110_0110_111: DATA = 1'b0;
            //VERTICAL LEFT 0 COL 0 Row 7
            15'b11000110_0111_000: DATA = 1'b1;
            15'b11000110_0111_001: DATA = 1'b0;
            15'b11000110_0111_010: DATA = 1'b0;
            15'b11000110_0111_011: DATA = 1'b0;
            15'b11000110_0111_100: DATA = 1'b0;
            15'b11000110_0111_101: DATA = 1'b0;
            15'b11000110_0111_110: DATA = 1'b0;
            15'b11000110_0111_111: DATA = 1'b0;
            //VERTICAL LEFT 0 COL 0 Row 8
            15'b11000110_1000_000: DATA = 1'b1;
            15'b11000110_1000_001: DATA = 1'b0;
            15'b11000110_1000_010: DATA = 1'b0;
            15'b11000110_1000_011: DATA = 1'b0;
            15'b11000110_1000_100: DATA = 1'b0;
            15'b11000110_1000_101: DATA = 1'b0;
            15'b11000110_1000_110: DATA = 1'b0;
            15'b11000110_1000_111: DATA = 1'b0;
            //VERTICAL LEFT 0 COL 0 Row 9
            15'b11000110_1001_000: DATA = 1'b1;
            15'b11000110_1001_001: DATA = 1'b0;
            15'b11000110_1001_010: DATA = 1'b0;
            15'b11000110_1001_011: DATA = 1'b0;
            15'b11000110_1001_100: DATA = 1'b0;
            15'b11000110_1001_101: DATA = 1'b0;
            15'b11000110_1001_110: DATA = 1'b0;
            15'b11000110_1001_111: DATA = 1'b0;
            //VERTICAL LEFT 0 COL 0 Row 10
            15'b11000110_1010_000: DATA = 1'b1;
            15'b11000110_1010_001: DATA = 1'b0;
            15'b11000110_1010_010: DATA = 1'b0;
            15'b11000110_1010_011: DATA = 1'b0;
            15'b11000110_1010_100: DATA = 1'b0;
            15'b11000110_1010_101: DATA = 1'b0;
            15'b11000110_1010_110: DATA = 1'b0;
            15'b11000110_1010_111: DATA = 1'b0;
            //VERTICAL LEFT 0 COL 0 Row 11
            15'b11000110_1011_000: DATA = 1'b1;
            15'b11000110_1011_001: DATA = 1'b0;
            15'b11000110_1011_010: DATA = 1'b0;
            15'b11000110_1011_011: DATA = 1'b0;
            15'b11000110_1011_100: DATA = 1'b0;
            15'b11000110_1011_101: DATA = 1'b0;
            15'b11000110_1011_110: DATA = 1'b0;
            15'b11000110_1011_111: DATA = 1'b0;
            //VERTICAL LEFT 0 COL 0 Row 12
            15'b11000110_1100_000: DATA = 1'b1;
            15'b11000110_1100_001: DATA = 1'b0;
            15'b11000110_1100_010: DATA = 1'b0;
            15'b11000110_1100_011: DATA = 1'b0;
            15'b11000110_1100_100: DATA = 1'b0;
            15'b11000110_1100_101: DATA = 1'b0;
            15'b11000110_1100_110: DATA = 1'b0;
            15'b11000110_1100_111: DATA = 1'b0;
            //VERTICAL LEFT 0 COL 0 Row 13
            15'b11000110_1101_000: DATA = 1'b1;
            15'b11000110_1101_001: DATA = 1'b0;
            15'b11000110_1101_010: DATA = 1'b0;
            15'b11000110_1101_011: DATA = 1'b0;
            15'b11000110_1101_100: DATA = 1'b0;
            15'b11000110_1101_101: DATA = 1'b0;
            15'b11000110_1101_110: DATA = 1'b0;
            15'b11000110_1101_111: DATA = 1'b0;
            //VERTICAL LEFT 0 COL 0 Row 14
            15'b11000110_1110_000: DATA = 1'b1;
            15'b11000110_1110_001: DATA = 1'b0;
            15'b11000110_1110_010: DATA = 1'b0;
            15'b11000110_1110_011: DATA = 1'b0;
            15'b11000110_1110_100: DATA = 1'b0;
            15'b11000110_1110_101: DATA = 1'b0;
            15'b11000110_1110_110: DATA = 1'b0;
            15'b11000110_1110_111: DATA = 1'b0;
            //VERTICAL LEFT 0 COL 0 Row 15
            15'b11000110_1111_000: DATA = 1'b1;
            15'b11000110_1111_001: DATA = 1'b0;
            15'b11000110_1111_010: DATA = 1'b0;
            15'b11000110_1111_011: DATA = 1'b0;
            15'b11000110_1111_100: DATA = 1'b0;
            15'b11000110_1111_101: DATA = 1'b0;
            15'b11000110_1111_110: DATA = 1'b0;
            15'b11000110_1111_111: DATA = 1'b0;
            //VERTICAL RIGHT 0 COL 0 Row 0
            15'b11000111_0000_000: DATA = 1'b0;
            15'b11000111_0000_001: DATA = 1'b0;
            15'b11000111_0000_010: DATA = 1'b0;
            15'b11000111_0000_011: DATA = 1'b0;
            15'b11000111_0000_100: DATA = 1'b0;
            15'b11000111_0000_101: DATA = 1'b0;
            15'b11000111_0000_110: DATA = 1'b0;
            15'b11000111_0000_111: DATA = 1'b1;
            //VERTICAL RIGHT 0 COL 0 Row 1
            15'b11000111_0001_000: DATA = 1'b0;
            15'b11000111_0001_001: DATA = 1'b0;
            15'b11000111_0001_010: DATA = 1'b0;
            15'b11000111_0001_011: DATA = 1'b0;
            15'b11000111_0001_100: DATA = 1'b0;
            15'b11000111_0001_101: DATA = 1'b0;
            15'b11000111_0001_110: DATA = 1'b0;
            15'b11000111_0001_111: DATA = 1'b1;
            //VERTICAL RIGHT 0 COL 0 Row 2
            15'b11000111_0010_000: DATA = 1'b0;
            15'b11000111_0010_001: DATA = 1'b0;
            15'b11000111_0010_010: DATA = 1'b0;
            15'b11000111_0010_011: DATA = 1'b0;
            15'b11000111_0010_100: DATA = 1'b0;
            15'b11000111_0010_101: DATA = 1'b0;
            15'b11000111_0010_110: DATA = 1'b0;
            15'b11000111_0010_111: DATA = 1'b1;
            //VERTICAL RIGHT 0 COL 0 Row 3
            15'b11000111_0011_000: DATA = 1'b0;
            15'b11000111_0011_001: DATA = 1'b0;
            15'b11000111_0011_010: DATA = 1'b0;
            15'b11000111_0011_011: DATA = 1'b0;
            15'b11000111_0011_100: DATA = 1'b0;
            15'b11000111_0011_101: DATA = 1'b0;
            15'b11000111_0011_110: DATA = 1'b0;
            15'b11000111_0011_111: DATA = 1'b1;
            //VERTICAL RIGHT 0 COL 0 Row 4
            15'b11000111_0100_000: DATA = 1'b0;
            15'b11000111_0100_001: DATA = 1'b0;
            15'b11000111_0100_010: DATA = 1'b0;
            15'b11000111_0100_011: DATA = 1'b0;
            15'b11000111_0100_100: DATA = 1'b0;
            15'b11000111_0100_101: DATA = 1'b0;
            15'b11000111_0100_110: DATA = 1'b0;
            15'b11000111_0100_111: DATA = 1'b1;
            //VERTICAL RIGHT 0 COL 0 Row 5
            15'b11000111_0101_000: DATA = 1'b0;
            15'b11000111_0101_001: DATA = 1'b0;
            15'b11000111_0101_010: DATA = 1'b0;
            15'b11000111_0101_011: DATA = 1'b0;
            15'b11000111_0101_100: DATA = 1'b0;
            15'b11000111_0101_101: DATA = 1'b0;
            15'b11000111_0101_110: DATA = 1'b0;
            15'b11000111_0101_111: DATA = 1'b1;
            //VERTICAL RIGHT 0 COL 0 Row 6
            15'b11000111_0110_000: DATA = 1'b0;
            15'b11000111_0110_001: DATA = 1'b0;
            15'b11000111_0110_010: DATA = 1'b0;
            15'b11000111_0110_011: DATA = 1'b0;
            15'b11000111_0110_100: DATA = 1'b0;
            15'b11000111_0110_101: DATA = 1'b0;
            15'b11000111_0110_110: DATA = 1'b0;
            15'b11000111_0110_111: DATA = 1'b1;
            //VERTICAL RIGHT 0 COL 0 Row 7
            15'b11000111_0111_000: DATA = 1'b0;
            15'b11000111_0111_001: DATA = 1'b0;
            15'b11000111_0111_010: DATA = 1'b0;
            15'b11000111_0111_011: DATA = 1'b0;
            15'b11000111_0111_100: DATA = 1'b0;
            15'b11000111_0111_101: DATA = 1'b0;
            15'b11000111_0111_110: DATA = 1'b0;
            15'b11000111_0111_111: DATA = 1'b1;
            //VERTICAL RIGHT 0 COL 0 Row 8
            15'b11000111_1000_000: DATA = 1'b0;
            15'b11000111_1000_001: DATA = 1'b0;
            15'b11000111_1000_010: DATA = 1'b0;
            15'b11000111_1000_011: DATA = 1'b0;
            15'b11000111_1000_100: DATA = 1'b0;
            15'b11000111_1000_101: DATA = 1'b0;
            15'b11000111_1000_110: DATA = 1'b0;
            15'b11000111_1000_111: DATA = 1'b1;
            //VERTICAL RIGHT 0 COL 0 Row 9
            15'b11000111_1001_000: DATA = 1'b0;
            15'b11000111_1001_001: DATA = 1'b0;
            15'b11000111_1001_010: DATA = 1'b0;
            15'b11000111_1001_011: DATA = 1'b0;
            15'b11000111_1001_100: DATA = 1'b0;
            15'b11000111_1001_101: DATA = 1'b0;
            15'b11000111_1001_110: DATA = 1'b0;
            15'b11000111_1001_111: DATA = 1'b1;
            //VERTICAL RIGHT 0 COL 0 Row 10
            15'b11000111_1010_000: DATA = 1'b0;
            15'b11000111_1010_001: DATA = 1'b0;
            15'b11000111_1010_010: DATA = 1'b0;
            15'b11000111_1010_011: DATA = 1'b0;
            15'b11000111_1010_100: DATA = 1'b0;
            15'b11000111_1010_101: DATA = 1'b0;
            15'b11000111_1010_110: DATA = 1'b0;
            15'b11000111_1010_111: DATA = 1'b1;
            //VERTICAL RIGHT 0 COL 0 Row 11
            15'b11000111_1011_000: DATA = 1'b0;
            15'b11000111_1011_001: DATA = 1'b0;
            15'b11000111_1011_010: DATA = 1'b0;
            15'b11000111_1011_011: DATA = 1'b0;
            15'b11000111_1011_100: DATA = 1'b0;
            15'b11000111_1011_101: DATA = 1'b0;
            15'b11000111_1011_110: DATA = 1'b0;
            15'b11000111_1011_111: DATA = 1'b1;
            //VERTICAL RIGHT 0 COL 0 Row 12
            15'b11000111_1100_000: DATA = 1'b0;
            15'b11000111_1100_001: DATA = 1'b0;
            15'b11000111_1100_010: DATA = 1'b0;
            15'b11000111_1100_011: DATA = 1'b0;
            15'b11000111_1100_100: DATA = 1'b0;
            15'b11000111_1100_101: DATA = 1'b0;
            15'b11000111_1100_110: DATA = 1'b0;
            15'b11000111_1100_111: DATA = 1'b1;
            //VERTICAL RIGHT 0 COL 0 Row 13
            15'b11000111_1101_000: DATA = 1'b0;
            15'b11000111_1101_001: DATA = 1'b0;
            15'b11000111_1101_010: DATA = 1'b0;
            15'b11000111_1101_011: DATA = 1'b0;
            15'b11000111_1101_100: DATA = 1'b0;
            15'b11000111_1101_101: DATA = 1'b0;
            15'b11000111_1101_110: DATA = 1'b0;
            15'b11000111_1101_111: DATA = 1'b1;
            //VERTICAL RIGHT 0 COL 0 Row 14
            15'b11000111_1110_000: DATA = 1'b0;
            15'b11000111_1110_001: DATA = 1'b0;
            15'b11000111_1110_010: DATA = 1'b0;
            15'b11000111_1110_011: DATA = 1'b0;
            15'b11000111_1110_100: DATA = 1'b0;
            15'b11000111_1110_101: DATA = 1'b0;
            15'b11000111_1110_110: DATA = 1'b0;
            15'b11000111_1110_111: DATA = 1'b1;
            //VERTICAL RIGHT 0 COL 0 Row 15
            15'b11000111_1111_000: DATA = 1'b0;
            15'b11000111_1111_001: DATA = 1'b0;
            15'b11000111_1111_010: DATA = 1'b0;
            15'b11000111_1111_011: DATA = 1'b0;
            15'b11000111_1111_100: DATA = 1'b0;
            15'b11000111_1111_101: DATA = 1'b0;
            15'b11000111_1111_110: DATA = 1'b0;
            15'b11000111_1111_111: DATA = 1'b1;
            //HORIZONTAL TOP 0 COL 0 Row 0
            15'b11001000_0000_000: DATA = 1'b1;
            15'b11001000_0000_001: DATA = 1'b1;
            15'b11001000_0000_010: DATA = 1'b1;
            15'b11001000_0000_011: DATA = 1'b1;
            15'b11001000_0000_100: DATA = 1'b1;
            15'b11001000_0000_101: DATA = 1'b1;
            15'b11001000_0000_110: DATA = 1'b1;
            15'b11001000_0000_111: DATA = 1'b1;
            //HORIZONTAL TOP 0 COL 0 Row 1
            15'b11001000_0001_000: DATA = 1'b0;
            15'b11001000_0001_001: DATA = 1'b0;
            15'b11001000_0001_010: DATA = 1'b0;
            15'b11001000_0001_011: DATA = 1'b0;
            15'b11001000_0001_100: DATA = 1'b0;
            15'b11001000_0001_101: DATA = 1'b0;
            15'b11001000_0001_110: DATA = 1'b0;
            15'b11001000_0001_111: DATA = 1'b0;
            //HORIZONTAL TOP 0 COL 0 Row 2
            15'b11001000_0010_000: DATA = 1'b0;
            15'b11001000_0010_001: DATA = 1'b0;
            15'b11001000_0010_010: DATA = 1'b0;
            15'b11001000_0010_011: DATA = 1'b0;
            15'b11001000_0010_100: DATA = 1'b0;
            15'b11001000_0010_101: DATA = 1'b0;
            15'b11001000_0010_110: DATA = 1'b0;
            15'b11001000_0010_111: DATA = 1'b0;
            //HORIZONTAL TOP 0 COL 0 Row 3
            15'b11001000_0011_000: DATA = 1'b0;
            15'b11001000_0011_001: DATA = 1'b0;
            15'b11001000_0011_010: DATA = 1'b0;
            15'b11001000_0011_011: DATA = 1'b0;
            15'b11001000_0011_100: DATA = 1'b0;
            15'b11001000_0011_101: DATA = 1'b0;
            15'b11001000_0011_110: DATA = 1'b0;
            15'b11001000_0011_111: DATA = 1'b0;
            //HORIZONTAL TOP 0 COL 0 Row 4
            15'b11001000_0100_000: DATA = 1'b0;
            15'b11001000_0100_001: DATA = 1'b0;
            15'b11001000_0100_010: DATA = 1'b0;
            15'b11001000_0100_011: DATA = 1'b0;
            15'b11001000_0100_100: DATA = 1'b0;
            15'b11001000_0100_101: DATA = 1'b0;
            15'b11001000_0100_110: DATA = 1'b0;
            15'b11001000_0100_111: DATA = 1'b0;
            //HORIZONTAL TOP 0 COL 0 Row 5
            15'b11001000_0101_000: DATA = 1'b0;
            15'b11001000_0101_001: DATA = 1'b0;
            15'b11001000_0101_010: DATA = 1'b0;
            15'b11001000_0101_011: DATA = 1'b0;
            15'b11001000_0101_100: DATA = 1'b0;
            15'b11001000_0101_101: DATA = 1'b0;
            15'b11001000_0101_110: DATA = 1'b0;
            15'b11001000_0101_111: DATA = 1'b0;
            //HORIZONTAL TOP 0 COL 0 Row 6
            15'b11001000_0110_000: DATA = 1'b0;
            15'b11001000_0110_001: DATA = 1'b0;
            15'b11001000_0110_010: DATA = 1'b0;
            15'b11001000_0110_011: DATA = 1'b0;
            15'b11001000_0110_100: DATA = 1'b0;
            15'b11001000_0110_101: DATA = 1'b0;
            15'b11001000_0110_110: DATA = 1'b0;
            15'b11001000_0110_111: DATA = 1'b0;
            //HORIZONTAL TOP 0 COL 0 Row 7
            15'b11001000_0111_000: DATA = 1'b0;
            15'b11001000_0111_001: DATA = 1'b0;
            15'b11001000_0111_010: DATA = 1'b0;
            15'b11001000_0111_011: DATA = 1'b0;
            15'b11001000_0111_100: DATA = 1'b0;
            15'b11001000_0111_101: DATA = 1'b0;
            15'b11001000_0111_110: DATA = 1'b0;
            15'b11001000_0111_111: DATA = 1'b0;
            //HORIZONTAL TOP 0 COL 0 Row 8
            15'b11001000_1000_000: DATA = 1'b0;
            15'b11001000_1000_001: DATA = 1'b0;
            15'b11001000_1000_010: DATA = 1'b0;
            15'b11001000_1000_011: DATA = 1'b0;
            15'b11001000_1000_100: DATA = 1'b0;
            15'b11001000_1000_101: DATA = 1'b0;
            15'b11001000_1000_110: DATA = 1'b0;
            15'b11001000_1000_111: DATA = 1'b0;
            //HORIZONTAL TOP 0 COL 0 Row 9
            15'b11001000_1001_000: DATA = 1'b0;
            15'b11001000_1001_001: DATA = 1'b0;
            15'b11001000_1001_010: DATA = 1'b0;
            15'b11001000_1001_011: DATA = 1'b0;
            15'b11001000_1001_100: DATA = 1'b0;
            15'b11001000_1001_101: DATA = 1'b0;
            15'b11001000_1001_110: DATA = 1'b0;
            15'b11001000_1001_111: DATA = 1'b0;
            //HORIZONTAL TOP 0 COL 0 Row 10
            15'b11001000_1010_000: DATA = 1'b0;
            15'b11001000_1010_001: DATA = 1'b0;
            15'b11001000_1010_010: DATA = 1'b0;
            15'b11001000_1010_011: DATA = 1'b0;
            15'b11001000_1010_100: DATA = 1'b0;
            15'b11001000_1010_101: DATA = 1'b0;
            15'b11001000_1010_110: DATA = 1'b0;
            15'b11001000_1010_111: DATA = 1'b0;
            //HORIZONTAL TOP 0 COL 0 Row 11
            15'b11001000_1011_000: DATA = 1'b0;
            15'b11001000_1011_001: DATA = 1'b0;
            15'b11001000_1011_010: DATA = 1'b0;
            15'b11001000_1011_011: DATA = 1'b0;
            15'b11001000_1011_100: DATA = 1'b0;
            15'b11001000_1011_101: DATA = 1'b0;
            15'b11001000_1011_110: DATA = 1'b0;
            15'b11001000_1011_111: DATA = 1'b0;
            //HORIZONTAL TOP 0 COL 0 Row 12
            15'b11001000_1100_000: DATA = 1'b0;
            15'b11001000_1100_001: DATA = 1'b0;
            15'b11001000_1100_010: DATA = 1'b0;
            15'b11001000_1100_011: DATA = 1'b0;
            15'b11001000_1100_100: DATA = 1'b0;
            15'b11001000_1100_101: DATA = 1'b0;
            15'b11001000_1100_110: DATA = 1'b0;
            15'b11001000_1100_111: DATA = 1'b0;
            //HORIZONTAL TOP 0 COL 0 Row 13
            15'b11001000_1101_000: DATA = 1'b0;
            15'b11001000_1101_001: DATA = 1'b0;
            15'b11001000_1101_010: DATA = 1'b0;
            15'b11001000_1101_011: DATA = 1'b0;
            15'b11001000_1101_100: DATA = 1'b0;
            15'b11001000_1101_101: DATA = 1'b0;
            15'b11001000_1101_110: DATA = 1'b0;
            15'b11001000_1101_111: DATA = 1'b0;
            //HORIZONTAL TOP 0 COL 0 Row 14
            15'b11001000_1110_000: DATA = 1'b0;
            15'b11001000_1110_001: DATA = 1'b0;
            15'b11001000_1110_010: DATA = 1'b0;
            15'b11001000_1110_011: DATA = 1'b0;
            15'b11001000_1110_100: DATA = 1'b0;
            15'b11001000_1110_101: DATA = 1'b0;
            15'b11001000_1110_110: DATA = 1'b0;
            15'b11001000_1110_111: DATA = 1'b0;
            //HORIZONTAL TOP 0 COL 0 Row 15
            15'b11001000_1111_000: DATA = 1'b0;
            15'b11001000_1111_001: DATA = 1'b0;
            15'b11001000_1111_010: DATA = 1'b0;
            15'b11001000_1111_011: DATA = 1'b0;
            15'b11001000_1111_100: DATA = 1'b0;
            15'b11001000_1111_101: DATA = 1'b0;
            15'b11001000_1111_110: DATA = 1'b0;
            15'b11001000_1111_111: DATA = 1'b0;
            //HORIZONTAL BOTTOM 0 COL 0 Row 0
            15'b11001001_0000_000: DATA = 1'b0;
            15'b11001001_0000_001: DATA = 1'b0;
            15'b11001001_0000_010: DATA = 1'b0;
            15'b11001001_0000_011: DATA = 1'b0;
            15'b11001001_0000_100: DATA = 1'b0;
            15'b11001001_0000_101: DATA = 1'b0;
            15'b11001001_0000_110: DATA = 1'b0;
            15'b11001001_0000_111: DATA = 1'b0;
            //HORIZONTAL BOTTOM 0 COL 0 Row 1
            15'b11001001_0001_000: DATA = 1'b0;
            15'b11001001_0001_001: DATA = 1'b0;
            15'b11001001_0001_010: DATA = 1'b0;
            15'b11001001_0001_011: DATA = 1'b0;
            15'b11001001_0001_100: DATA = 1'b0;
            15'b11001001_0001_101: DATA = 1'b0;
            15'b11001001_0001_110: DATA = 1'b0;
            15'b11001001_0001_111: DATA = 1'b0;
            //HORIZONTAL BOTTOM 0 COL 0 Row 2
            15'b11001001_0010_000: DATA = 1'b0;
            15'b11001001_0010_001: DATA = 1'b0;
            15'b11001001_0010_010: DATA = 1'b0;
            15'b11001001_0010_011: DATA = 1'b0;
            15'b11001001_0010_100: DATA = 1'b0;
            15'b11001001_0010_101: DATA = 1'b0;
            15'b11001001_0010_110: DATA = 1'b0;
            15'b11001001_0010_111: DATA = 1'b0;
            //HORIZONTAL BOTTOM 0 COL 0 Row 3
            15'b11001001_0011_000: DATA = 1'b0;
            15'b11001001_0011_001: DATA = 1'b0;
            15'b11001001_0011_010: DATA = 1'b0;
            15'b11001001_0011_011: DATA = 1'b0;
            15'b11001001_0011_100: DATA = 1'b0;
            15'b11001001_0011_101: DATA = 1'b0;
            15'b11001001_0011_110: DATA = 1'b0;
            15'b11001001_0011_111: DATA = 1'b0;
            //HORIZONTAL BOTTOM 0 COL 0 Row 4
            15'b11001001_0100_000: DATA = 1'b0;
            15'b11001001_0100_001: DATA = 1'b0;
            15'b11001001_0100_010: DATA = 1'b0;
            15'b11001001_0100_011: DATA = 1'b0;
            15'b11001001_0100_100: DATA = 1'b0;
            15'b11001001_0100_101: DATA = 1'b0;
            15'b11001001_0100_110: DATA = 1'b0;
            15'b11001001_0100_111: DATA = 1'b0;
            //HORIZONTAL BOTTOM 0 COL 0 Row 5
            15'b11001001_0101_000: DATA = 1'b0;
            15'b11001001_0101_001: DATA = 1'b0;
            15'b11001001_0101_010: DATA = 1'b0;
            15'b11001001_0101_011: DATA = 1'b0;
            15'b11001001_0101_100: DATA = 1'b0;
            15'b11001001_0101_101: DATA = 1'b0;
            15'b11001001_0101_110: DATA = 1'b0;
            15'b11001001_0101_111: DATA = 1'b0;
            //HORIZONTAL BOTTOM 0 COL 0 Row 6
            15'b11001001_0110_000: DATA = 1'b0;
            15'b11001001_0110_001: DATA = 1'b0;
            15'b11001001_0110_010: DATA = 1'b0;
            15'b11001001_0110_011: DATA = 1'b0;
            15'b11001001_0110_100: DATA = 1'b0;
            15'b11001001_0110_101: DATA = 1'b0;
            15'b11001001_0110_110: DATA = 1'b0;
            15'b11001001_0110_111: DATA = 1'b0;
            //HORIZONTAL BOTTOM 0 COL 0 Row 7
            15'b11001001_0111_000: DATA = 1'b0;
            15'b11001001_0111_001: DATA = 1'b0;
            15'b11001001_0111_010: DATA = 1'b0;
            15'b11001001_0111_011: DATA = 1'b0;
            15'b11001001_0111_100: DATA = 1'b0;
            15'b11001001_0111_101: DATA = 1'b0;
            15'b11001001_0111_110: DATA = 1'b0;
            15'b11001001_0111_111: DATA = 1'b0;
            //HORIZONTAL BOTTOM 0 COL 0 Row 8
            15'b11001001_1000_000: DATA = 1'b0;
            15'b11001001_1000_001: DATA = 1'b0;
            15'b11001001_1000_010: DATA = 1'b0;
            15'b11001001_1000_011: DATA = 1'b0;
            15'b11001001_1000_100: DATA = 1'b0;
            15'b11001001_1000_101: DATA = 1'b0;
            15'b11001001_1000_110: DATA = 1'b0;
            15'b11001001_1000_111: DATA = 1'b0;
            //HORIZONTAL BOTTOM 0 COL 0 Row 9
            15'b11001001_1001_000: DATA = 1'b0;
            15'b11001001_1001_001: DATA = 1'b0;
            15'b11001001_1001_010: DATA = 1'b0;
            15'b11001001_1001_011: DATA = 1'b0;
            15'b11001001_1001_100: DATA = 1'b0;
            15'b11001001_1001_101: DATA = 1'b0;
            15'b11001001_1001_110: DATA = 1'b0;
            15'b11001001_1001_111: DATA = 1'b0;
            //HORIZONTAL BOTTOM 0 COL 0 Row 10
            15'b11001001_1010_000: DATA = 1'b0;
            15'b11001001_1010_001: DATA = 1'b0;
            15'b11001001_1010_010: DATA = 1'b0;
            15'b11001001_1010_011: DATA = 1'b0;
            15'b11001001_1010_100: DATA = 1'b0;
            15'b11001001_1010_101: DATA = 1'b0;
            15'b11001001_1010_110: DATA = 1'b0;
            15'b11001001_1010_111: DATA = 1'b0;
            //HORIZONTAL BOTTOM 0 COL 0 Row 11
            15'b11001001_1011_000: DATA = 1'b0;
            15'b11001001_1011_001: DATA = 1'b0;
            15'b11001001_1011_010: DATA = 1'b0;
            15'b11001001_1011_011: DATA = 1'b0;
            15'b11001001_1011_100: DATA = 1'b0;
            15'b11001001_1011_101: DATA = 1'b0;
            15'b11001001_1011_110: DATA = 1'b0;
            15'b11001001_1011_111: DATA = 1'b0;
            //HORIZONTAL BOTTOM 0 COL 0 Row 12
            15'b11001001_1100_000: DATA = 1'b0;
            15'b11001001_1100_001: DATA = 1'b0;
            15'b11001001_1100_010: DATA = 1'b0;
            15'b11001001_1100_011: DATA = 1'b0;
            15'b11001001_1100_100: DATA = 1'b0;
            15'b11001001_1100_101: DATA = 1'b0;
            15'b11001001_1100_110: DATA = 1'b0;
            15'b11001001_1100_111: DATA = 1'b0;
            //HORIZONTAL BOTTOM 0 COL 0 Row 13
            15'b11001001_1101_000: DATA = 1'b0;
            15'b11001001_1101_001: DATA = 1'b0;
            15'b11001001_1101_010: DATA = 1'b0;
            15'b11001001_1101_011: DATA = 1'b0;
            15'b11001001_1101_100: DATA = 1'b0;
            15'b11001001_1101_101: DATA = 1'b0;
            15'b11001001_1101_110: DATA = 1'b0;
            15'b11001001_1101_111: DATA = 1'b0;
            //HORIZONTAL BOTTOM 0 COL 0 Row 14
            15'b11001001_1110_000: DATA = 1'b0;
            15'b11001001_1110_001: DATA = 1'b0;
            15'b11001001_1110_010: DATA = 1'b0;
            15'b11001001_1110_011: DATA = 1'b0;
            15'b11001001_1110_100: DATA = 1'b0;
            15'b11001001_1110_101: DATA = 1'b0;
            15'b11001001_1110_110: DATA = 1'b0;
            15'b11001001_1110_111: DATA = 1'b0;
            //HORIZONTAL BOTTOM 0 COL 0 Row 15
            15'b11001001_1111_000: DATA = 1'b1;
            15'b11001001_1111_001: DATA = 1'b1;
            15'b11001001_1111_010: DATA = 1'b1;
            15'b11001001_1111_011: DATA = 1'b1;
            15'b11001001_1111_100: DATA = 1'b1;
            15'b11001001_1111_101: DATA = 1'b1;
            15'b11001001_1111_110: DATA = 1'b1;
            15'b11001001_1111_111: DATA = 1'b1;
            //SAWTOOTH- ROW 0 COL 0 Row 0
            15'b11001010_0000_000: DATA = 1'b1;
            15'b11001010_0000_001: DATA = 1'b0;
            15'b11001010_0000_010: DATA = 1'b0;
            15'b11001010_0000_011: DATA = 1'b0;
            15'b11001010_0000_100: DATA = 1'b0;
            15'b11001010_0000_101: DATA = 1'b0;
            15'b11001010_0000_110: DATA = 1'b0;
            15'b11001010_0000_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 0 Row 1
            15'b11001010_0001_000: DATA = 1'b1;
            15'b11001010_0001_001: DATA = 1'b0;
            15'b11001010_0001_010: DATA = 1'b0;
            15'b11001010_0001_011: DATA = 1'b0;
            15'b11001010_0001_100: DATA = 1'b0;
            15'b11001010_0001_101: DATA = 1'b0;
            15'b11001010_0001_110: DATA = 1'b0;
            15'b11001010_0001_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 0 Row 2
            15'b11001010_0010_000: DATA = 1'b1;
            15'b11001010_0010_001: DATA = 1'b0;
            15'b11001010_0010_010: DATA = 1'b0;
            15'b11001010_0010_011: DATA = 1'b0;
            15'b11001010_0010_100: DATA = 1'b0;
            15'b11001010_0010_101: DATA = 1'b0;
            15'b11001010_0010_110: DATA = 1'b0;
            15'b11001010_0010_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 0 Row 3
            15'b11001010_0011_000: DATA = 1'b1;
            15'b11001010_0011_001: DATA = 1'b0;
            15'b11001010_0011_010: DATA = 1'b0;
            15'b11001010_0011_011: DATA = 1'b0;
            15'b11001010_0011_100: DATA = 1'b0;
            15'b11001010_0011_101: DATA = 1'b0;
            15'b11001010_0011_110: DATA = 1'b0;
            15'b11001010_0011_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 0 Row 4
            15'b11001010_0100_000: DATA = 1'b1;
            15'b11001010_0100_001: DATA = 1'b0;
            15'b11001010_0100_010: DATA = 1'b0;
            15'b11001010_0100_011: DATA = 1'b0;
            15'b11001010_0100_100: DATA = 1'b0;
            15'b11001010_0100_101: DATA = 1'b0;
            15'b11001010_0100_110: DATA = 1'b0;
            15'b11001010_0100_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 0 Row 5
            15'b11001010_0101_000: DATA = 1'b1;
            15'b11001010_0101_001: DATA = 1'b0;
            15'b11001010_0101_010: DATA = 1'b0;
            15'b11001010_0101_011: DATA = 1'b0;
            15'b11001010_0101_100: DATA = 1'b0;
            15'b11001010_0101_101: DATA = 1'b0;
            15'b11001010_0101_110: DATA = 1'b0;
            15'b11001010_0101_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 0 Row 6
            15'b11001010_0110_000: DATA = 1'b1;
            15'b11001010_0110_001: DATA = 1'b0;
            15'b11001010_0110_010: DATA = 1'b0;
            15'b11001010_0110_011: DATA = 1'b0;
            15'b11001010_0110_100: DATA = 1'b0;
            15'b11001010_0110_101: DATA = 1'b0;
            15'b11001010_0110_110: DATA = 1'b0;
            15'b11001010_0110_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 0 Row 7
            15'b11001010_0111_000: DATA = 1'b1;
            15'b11001010_0111_001: DATA = 1'b0;
            15'b11001010_0111_010: DATA = 1'b0;
            15'b11001010_0111_011: DATA = 1'b0;
            15'b11001010_0111_100: DATA = 1'b0;
            15'b11001010_0111_101: DATA = 1'b0;
            15'b11001010_0111_110: DATA = 1'b0;
            15'b11001010_0111_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 0 Row 8
            15'b11001010_1000_000: DATA = 1'b1;
            15'b11001010_1000_001: DATA = 1'b0;
            15'b11001010_1000_010: DATA = 1'b0;
            15'b11001010_1000_011: DATA = 1'b0;
            15'b11001010_1000_100: DATA = 1'b0;
            15'b11001010_1000_101: DATA = 1'b0;
            15'b11001010_1000_110: DATA = 1'b0;
            15'b11001010_1000_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 0 Row 9
            15'b11001010_1001_000: DATA = 1'b1;
            15'b11001010_1001_001: DATA = 1'b0;
            15'b11001010_1001_010: DATA = 1'b0;
            15'b11001010_1001_011: DATA = 1'b0;
            15'b11001010_1001_100: DATA = 1'b0;
            15'b11001010_1001_101: DATA = 1'b0;
            15'b11001010_1001_110: DATA = 1'b0;
            15'b11001010_1001_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 0 Row 10
            15'b11001010_1010_000: DATA = 1'b1;
            15'b11001010_1010_001: DATA = 1'b0;
            15'b11001010_1010_010: DATA = 1'b0;
            15'b11001010_1010_011: DATA = 1'b0;
            15'b11001010_1010_100: DATA = 1'b0;
            15'b11001010_1010_101: DATA = 1'b0;
            15'b11001010_1010_110: DATA = 1'b0;
            15'b11001010_1010_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 0 Row 11
            15'b11001010_1011_000: DATA = 1'b1;
            15'b11001010_1011_001: DATA = 1'b0;
            15'b11001010_1011_010: DATA = 1'b0;
            15'b11001010_1011_011: DATA = 1'b0;
            15'b11001010_1011_100: DATA = 1'b0;
            15'b11001010_1011_101: DATA = 1'b0;
            15'b11001010_1011_110: DATA = 1'b0;
            15'b11001010_1011_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 0 Row 12
            15'b11001010_1100_000: DATA = 1'b1;
            15'b11001010_1100_001: DATA = 1'b0;
            15'b11001010_1100_010: DATA = 1'b0;
            15'b11001010_1100_011: DATA = 1'b0;
            15'b11001010_1100_100: DATA = 1'b0;
            15'b11001010_1100_101: DATA = 1'b0;
            15'b11001010_1100_110: DATA = 1'b0;
            15'b11001010_1100_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 0 Row 13
            15'b11001010_1101_000: DATA = 1'b1;
            15'b11001010_1101_001: DATA = 1'b0;
            15'b11001010_1101_010: DATA = 1'b0;
            15'b11001010_1101_011: DATA = 1'b0;
            15'b11001010_1101_100: DATA = 1'b0;
            15'b11001010_1101_101: DATA = 1'b0;
            15'b11001010_1101_110: DATA = 1'b0;
            15'b11001010_1101_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 0 Row 14
            15'b11001010_1110_000: DATA = 1'b1;
            15'b11001010_1110_001: DATA = 1'b0;
            15'b11001010_1110_010: DATA = 1'b0;
            15'b11001010_1110_011: DATA = 1'b0;
            15'b11001010_1110_100: DATA = 1'b0;
            15'b11001010_1110_101: DATA = 1'b0;
            15'b11001010_1110_110: DATA = 1'b0;
            15'b11001010_1110_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 0 Row 15
            15'b11001010_1111_000: DATA = 1'b1;
            15'b11001010_1111_001: DATA = 1'b0;
            15'b11001010_1111_010: DATA = 1'b0;
            15'b11001010_1111_011: DATA = 1'b0;
            15'b11001010_1111_100: DATA = 1'b0;
            15'b11001010_1111_101: DATA = 1'b0;
            15'b11001010_1111_110: DATA = 1'b0;
            15'b11001010_1111_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 1 Row 0
            15'b11001011_0000_000: DATA = 1'b0;
            15'b11001011_0000_001: DATA = 1'b0;
            15'b11001011_0000_010: DATA = 1'b0;
            15'b11001011_0000_011: DATA = 1'b0;
            15'b11001011_0000_100: DATA = 1'b0;
            15'b11001011_0000_101: DATA = 1'b0;
            15'b11001011_0000_110: DATA = 1'b0;
            15'b11001011_0000_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 1 Row 1
            15'b11001011_0001_000: DATA = 1'b0;
            15'b11001011_0001_001: DATA = 1'b0;
            15'b11001011_0001_010: DATA = 1'b0;
            15'b11001011_0001_011: DATA = 1'b0;
            15'b11001011_0001_100: DATA = 1'b0;
            15'b11001011_0001_101: DATA = 1'b0;
            15'b11001011_0001_110: DATA = 1'b0;
            15'b11001011_0001_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 1 Row 2
            15'b11001011_0010_000: DATA = 1'b0;
            15'b11001011_0010_001: DATA = 1'b0;
            15'b11001011_0010_010: DATA = 1'b0;
            15'b11001011_0010_011: DATA = 1'b0;
            15'b11001011_0010_100: DATA = 1'b0;
            15'b11001011_0010_101: DATA = 1'b0;
            15'b11001011_0010_110: DATA = 1'b0;
            15'b11001011_0010_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 1 Row 3
            15'b11001011_0011_000: DATA = 1'b0;
            15'b11001011_0011_001: DATA = 1'b0;
            15'b11001011_0011_010: DATA = 1'b0;
            15'b11001011_0011_011: DATA = 1'b0;
            15'b11001011_0011_100: DATA = 1'b0;
            15'b11001011_0011_101: DATA = 1'b0;
            15'b11001011_0011_110: DATA = 1'b0;
            15'b11001011_0011_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 1 Row 4
            15'b11001011_0100_000: DATA = 1'b0;
            15'b11001011_0100_001: DATA = 1'b0;
            15'b11001011_0100_010: DATA = 1'b0;
            15'b11001011_0100_011: DATA = 1'b0;
            15'b11001011_0100_100: DATA = 1'b0;
            15'b11001011_0100_101: DATA = 1'b0;
            15'b11001011_0100_110: DATA = 1'b0;
            15'b11001011_0100_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 1 Row 5
            15'b11001011_0101_000: DATA = 1'b0;
            15'b11001011_0101_001: DATA = 1'b0;
            15'b11001011_0101_010: DATA = 1'b0;
            15'b11001011_0101_011: DATA = 1'b0;
            15'b11001011_0101_100: DATA = 1'b0;
            15'b11001011_0101_101: DATA = 1'b0;
            15'b11001011_0101_110: DATA = 1'b0;
            15'b11001011_0101_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 1 Row 6
            15'b11001011_0110_000: DATA = 1'b0;
            15'b11001011_0110_001: DATA = 1'b0;
            15'b11001011_0110_010: DATA = 1'b0;
            15'b11001011_0110_011: DATA = 1'b0;
            15'b11001011_0110_100: DATA = 1'b0;
            15'b11001011_0110_101: DATA = 1'b0;
            15'b11001011_0110_110: DATA = 1'b0;
            15'b11001011_0110_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 1 Row 7
            15'b11001011_0111_000: DATA = 1'b0;
            15'b11001011_0111_001: DATA = 1'b0;
            15'b11001011_0111_010: DATA = 1'b0;
            15'b11001011_0111_011: DATA = 1'b0;
            15'b11001011_0111_100: DATA = 1'b0;
            15'b11001011_0111_101: DATA = 1'b0;
            15'b11001011_0111_110: DATA = 1'b0;
            15'b11001011_0111_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 1 Row 8
            15'b11001011_1000_000: DATA = 1'b0;
            15'b11001011_1000_001: DATA = 1'b0;
            15'b11001011_1000_010: DATA = 1'b0;
            15'b11001011_1000_011: DATA = 1'b0;
            15'b11001011_1000_100: DATA = 1'b0;
            15'b11001011_1000_101: DATA = 1'b0;
            15'b11001011_1000_110: DATA = 1'b0;
            15'b11001011_1000_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 1 Row 9
            15'b11001011_1001_000: DATA = 1'b0;
            15'b11001011_1001_001: DATA = 1'b0;
            15'b11001011_1001_010: DATA = 1'b0;
            15'b11001011_1001_011: DATA = 1'b0;
            15'b11001011_1001_100: DATA = 1'b0;
            15'b11001011_1001_101: DATA = 1'b0;
            15'b11001011_1001_110: DATA = 1'b0;
            15'b11001011_1001_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 1 Row 10
            15'b11001011_1010_000: DATA = 1'b0;
            15'b11001011_1010_001: DATA = 1'b0;
            15'b11001011_1010_010: DATA = 1'b0;
            15'b11001011_1010_011: DATA = 1'b0;
            15'b11001011_1010_100: DATA = 1'b0;
            15'b11001011_1010_101: DATA = 1'b0;
            15'b11001011_1010_110: DATA = 1'b0;
            15'b11001011_1010_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 1 Row 11
            15'b11001011_1011_000: DATA = 1'b0;
            15'b11001011_1011_001: DATA = 1'b0;
            15'b11001011_1011_010: DATA = 1'b0;
            15'b11001011_1011_011: DATA = 1'b0;
            15'b11001011_1011_100: DATA = 1'b0;
            15'b11001011_1011_101: DATA = 1'b0;
            15'b11001011_1011_110: DATA = 1'b0;
            15'b11001011_1011_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 1 Row 12
            15'b11001011_1100_000: DATA = 1'b0;
            15'b11001011_1100_001: DATA = 1'b0;
            15'b11001011_1100_010: DATA = 1'b0;
            15'b11001011_1100_011: DATA = 1'b0;
            15'b11001011_1100_100: DATA = 1'b0;
            15'b11001011_1100_101: DATA = 1'b0;
            15'b11001011_1100_110: DATA = 1'b0;
            15'b11001011_1100_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 1 Row 13
            15'b11001011_1101_000: DATA = 1'b0;
            15'b11001011_1101_001: DATA = 1'b0;
            15'b11001011_1101_010: DATA = 1'b0;
            15'b11001011_1101_011: DATA = 1'b0;
            15'b11001011_1101_100: DATA = 1'b0;
            15'b11001011_1101_101: DATA = 1'b0;
            15'b11001011_1101_110: DATA = 1'b0;
            15'b11001011_1101_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 1 Row 14
            15'b11001011_1110_000: DATA = 1'b0;
            15'b11001011_1110_001: DATA = 1'b0;
            15'b11001011_1110_010: DATA = 1'b0;
            15'b11001011_1110_011: DATA = 1'b0;
            15'b11001011_1110_100: DATA = 1'b0;
            15'b11001011_1110_101: DATA = 1'b0;
            15'b11001011_1110_110: DATA = 1'b0;
            15'b11001011_1110_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 1 Row 15
            15'b11001011_1111_000: DATA = 1'b0;
            15'b11001011_1111_001: DATA = 1'b0;
            15'b11001011_1111_010: DATA = 1'b0;
            15'b11001011_1111_011: DATA = 1'b0;
            15'b11001011_1111_100: DATA = 1'b0;
            15'b11001011_1111_101: DATA = 1'b0;
            15'b11001011_1111_110: DATA = 1'b0;
            15'b11001011_1111_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 2 Row 0
            15'b11001100_0000_000: DATA = 1'b0;
            15'b11001100_0000_001: DATA = 1'b0;
            15'b11001100_0000_010: DATA = 1'b0;
            15'b11001100_0000_011: DATA = 1'b0;
            15'b11001100_0000_100: DATA = 1'b0;
            15'b11001100_0000_101: DATA = 1'b0;
            15'b11001100_0000_110: DATA = 1'b0;
            15'b11001100_0000_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 2 Row 1
            15'b11001100_0001_000: DATA = 1'b0;
            15'b11001100_0001_001: DATA = 1'b0;
            15'b11001100_0001_010: DATA = 1'b0;
            15'b11001100_0001_011: DATA = 1'b0;
            15'b11001100_0001_100: DATA = 1'b0;
            15'b11001100_0001_101: DATA = 1'b0;
            15'b11001100_0001_110: DATA = 1'b0;
            15'b11001100_0001_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 2 Row 2
            15'b11001100_0010_000: DATA = 1'b0;
            15'b11001100_0010_001: DATA = 1'b0;
            15'b11001100_0010_010: DATA = 1'b0;
            15'b11001100_0010_011: DATA = 1'b0;
            15'b11001100_0010_100: DATA = 1'b0;
            15'b11001100_0010_101: DATA = 1'b0;
            15'b11001100_0010_110: DATA = 1'b0;
            15'b11001100_0010_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 2 Row 3
            15'b11001100_0011_000: DATA = 1'b0;
            15'b11001100_0011_001: DATA = 1'b0;
            15'b11001100_0011_010: DATA = 1'b0;
            15'b11001100_0011_011: DATA = 1'b0;
            15'b11001100_0011_100: DATA = 1'b0;
            15'b11001100_0011_101: DATA = 1'b0;
            15'b11001100_0011_110: DATA = 1'b0;
            15'b11001100_0011_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 2 Row 4
            15'b11001100_0100_000: DATA = 1'b0;
            15'b11001100_0100_001: DATA = 1'b0;
            15'b11001100_0100_010: DATA = 1'b0;
            15'b11001100_0100_011: DATA = 1'b0;
            15'b11001100_0100_100: DATA = 1'b0;
            15'b11001100_0100_101: DATA = 1'b0;
            15'b11001100_0100_110: DATA = 1'b0;
            15'b11001100_0100_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 2 Row 5
            15'b11001100_0101_000: DATA = 1'b0;
            15'b11001100_0101_001: DATA = 1'b0;
            15'b11001100_0101_010: DATA = 1'b0;
            15'b11001100_0101_011: DATA = 1'b0;
            15'b11001100_0101_100: DATA = 1'b0;
            15'b11001100_0101_101: DATA = 1'b0;
            15'b11001100_0101_110: DATA = 1'b0;
            15'b11001100_0101_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 2 Row 6
            15'b11001100_0110_000: DATA = 1'b0;
            15'b11001100_0110_001: DATA = 1'b0;
            15'b11001100_0110_010: DATA = 1'b0;
            15'b11001100_0110_011: DATA = 1'b0;
            15'b11001100_0110_100: DATA = 1'b0;
            15'b11001100_0110_101: DATA = 1'b0;
            15'b11001100_0110_110: DATA = 1'b0;
            15'b11001100_0110_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 2 Row 7
            15'b11001100_0111_000: DATA = 1'b0;
            15'b11001100_0111_001: DATA = 1'b0;
            15'b11001100_0111_010: DATA = 1'b0;
            15'b11001100_0111_011: DATA = 1'b0;
            15'b11001100_0111_100: DATA = 1'b0;
            15'b11001100_0111_101: DATA = 1'b0;
            15'b11001100_0111_110: DATA = 1'b0;
            15'b11001100_0111_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 2 Row 8
            15'b11001100_1000_000: DATA = 1'b0;
            15'b11001100_1000_001: DATA = 1'b0;
            15'b11001100_1000_010: DATA = 1'b0;
            15'b11001100_1000_011: DATA = 1'b0;
            15'b11001100_1000_100: DATA = 1'b0;
            15'b11001100_1000_101: DATA = 1'b0;
            15'b11001100_1000_110: DATA = 1'b0;
            15'b11001100_1000_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 2 Row 9
            15'b11001100_1001_000: DATA = 1'b0;
            15'b11001100_1001_001: DATA = 1'b0;
            15'b11001100_1001_010: DATA = 1'b0;
            15'b11001100_1001_011: DATA = 1'b0;
            15'b11001100_1001_100: DATA = 1'b0;
            15'b11001100_1001_101: DATA = 1'b0;
            15'b11001100_1001_110: DATA = 1'b0;
            15'b11001100_1001_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 2 Row 10
            15'b11001100_1010_000: DATA = 1'b0;
            15'b11001100_1010_001: DATA = 1'b0;
            15'b11001100_1010_010: DATA = 1'b0;
            15'b11001100_1010_011: DATA = 1'b0;
            15'b11001100_1010_100: DATA = 1'b0;
            15'b11001100_1010_101: DATA = 1'b0;
            15'b11001100_1010_110: DATA = 1'b0;
            15'b11001100_1010_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 2 Row 11
            15'b11001100_1011_000: DATA = 1'b0;
            15'b11001100_1011_001: DATA = 1'b0;
            15'b11001100_1011_010: DATA = 1'b0;
            15'b11001100_1011_011: DATA = 1'b0;
            15'b11001100_1011_100: DATA = 1'b0;
            15'b11001100_1011_101: DATA = 1'b0;
            15'b11001100_1011_110: DATA = 1'b0;
            15'b11001100_1011_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 2 Row 12
            15'b11001100_1100_000: DATA = 1'b0;
            15'b11001100_1100_001: DATA = 1'b0;
            15'b11001100_1100_010: DATA = 1'b0;
            15'b11001100_1100_011: DATA = 1'b0;
            15'b11001100_1100_100: DATA = 1'b0;
            15'b11001100_1100_101: DATA = 1'b0;
            15'b11001100_1100_110: DATA = 1'b0;
            15'b11001100_1100_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 2 Row 13
            15'b11001100_1101_000: DATA = 1'b0;
            15'b11001100_1101_001: DATA = 1'b0;
            15'b11001100_1101_010: DATA = 1'b0;
            15'b11001100_1101_011: DATA = 1'b0;
            15'b11001100_1101_100: DATA = 1'b0;
            15'b11001100_1101_101: DATA = 1'b0;
            15'b11001100_1101_110: DATA = 1'b0;
            15'b11001100_1101_111: DATA = 1'b1;
            //SAWTOOTH- ROW 0 COL 2 Row 14
            15'b11001100_1110_000: DATA = 1'b0;
            15'b11001100_1110_001: DATA = 1'b0;
            15'b11001100_1110_010: DATA = 1'b0;
            15'b11001100_1110_011: DATA = 1'b0;
            15'b11001100_1110_100: DATA = 1'b0;
            15'b11001100_1110_101: DATA = 1'b0;
            15'b11001100_1110_110: DATA = 1'b1;
            15'b11001100_1110_111: DATA = 1'b1;
            //SAWTOOTH- ROW 0 COL 2 Row 15
            15'b11001100_1111_000: DATA = 1'b0;
            15'b11001100_1111_001: DATA = 1'b0;
            15'b11001100_1111_010: DATA = 1'b0;
            15'b11001100_1111_011: DATA = 1'b0;
            15'b11001100_1111_100: DATA = 1'b0;
            15'b11001100_1111_101: DATA = 1'b1;
            15'b11001100_1111_110: DATA = 1'b1;
            15'b11001100_1111_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 3 Row 0
            15'b11001101_0000_000: DATA = 1'b0;
            15'b11001101_0000_001: DATA = 1'b0;
            15'b11001101_0000_010: DATA = 1'b0;
            15'b11001101_0000_011: DATA = 1'b0;
            15'b11001101_0000_100: DATA = 1'b0;
            15'b11001101_0000_101: DATA = 1'b0;
            15'b11001101_0000_110: DATA = 1'b0;
            15'b11001101_0000_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 3 Row 1
            15'b11001101_0001_000: DATA = 1'b0;
            15'b11001101_0001_001: DATA = 1'b0;
            15'b11001101_0001_010: DATA = 1'b0;
            15'b11001101_0001_011: DATA = 1'b0;
            15'b11001101_0001_100: DATA = 1'b0;
            15'b11001101_0001_101: DATA = 1'b0;
            15'b11001101_0001_110: DATA = 1'b0;
            15'b11001101_0001_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 3 Row 2
            15'b11001101_0010_000: DATA = 1'b0;
            15'b11001101_0010_001: DATA = 1'b0;
            15'b11001101_0010_010: DATA = 1'b0;
            15'b11001101_0010_011: DATA = 1'b0;
            15'b11001101_0010_100: DATA = 1'b0;
            15'b11001101_0010_101: DATA = 1'b0;
            15'b11001101_0010_110: DATA = 1'b0;
            15'b11001101_0010_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 3 Row 3
            15'b11001101_0011_000: DATA = 1'b0;
            15'b11001101_0011_001: DATA = 1'b0;
            15'b11001101_0011_010: DATA = 1'b0;
            15'b11001101_0011_011: DATA = 1'b0;
            15'b11001101_0011_100: DATA = 1'b0;
            15'b11001101_0011_101: DATA = 1'b0;
            15'b11001101_0011_110: DATA = 1'b0;
            15'b11001101_0011_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 3 Row 4
            15'b11001101_0100_000: DATA = 1'b0;
            15'b11001101_0100_001: DATA = 1'b0;
            15'b11001101_0100_010: DATA = 1'b0;
            15'b11001101_0100_011: DATA = 1'b0;
            15'b11001101_0100_100: DATA = 1'b0;
            15'b11001101_0100_101: DATA = 1'b0;
            15'b11001101_0100_110: DATA = 1'b0;
            15'b11001101_0100_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 3 Row 5
            15'b11001101_0101_000: DATA = 1'b0;
            15'b11001101_0101_001: DATA = 1'b0;
            15'b11001101_0101_010: DATA = 1'b0;
            15'b11001101_0101_011: DATA = 1'b0;
            15'b11001101_0101_100: DATA = 1'b0;
            15'b11001101_0101_101: DATA = 1'b0;
            15'b11001101_0101_110: DATA = 1'b0;
            15'b11001101_0101_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 3 Row 6
            15'b11001101_0110_000: DATA = 1'b0;
            15'b11001101_0110_001: DATA = 1'b0;
            15'b11001101_0110_010: DATA = 1'b0;
            15'b11001101_0110_011: DATA = 1'b0;
            15'b11001101_0110_100: DATA = 1'b0;
            15'b11001101_0110_101: DATA = 1'b0;
            15'b11001101_0110_110: DATA = 1'b0;
            15'b11001101_0110_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 3 Row 7
            15'b11001101_0111_000: DATA = 1'b0;
            15'b11001101_0111_001: DATA = 1'b0;
            15'b11001101_0111_010: DATA = 1'b0;
            15'b11001101_0111_011: DATA = 1'b0;
            15'b11001101_0111_100: DATA = 1'b0;
            15'b11001101_0111_101: DATA = 1'b0;
            15'b11001101_0111_110: DATA = 1'b0;
            15'b11001101_0111_111: DATA = 1'b1;
            //SAWTOOTH- ROW 0 COL 3 Row 8
            15'b11001101_1000_000: DATA = 1'b0;
            15'b11001101_1000_001: DATA = 1'b0;
            15'b11001101_1000_010: DATA = 1'b0;
            15'b11001101_1000_011: DATA = 1'b0;
            15'b11001101_1000_100: DATA = 1'b0;
            15'b11001101_1000_101: DATA = 1'b1;
            15'b11001101_1000_110: DATA = 1'b1;
            15'b11001101_1000_111: DATA = 1'b1;
            //SAWTOOTH- ROW 0 COL 3 Row 9
            15'b11001101_1001_000: DATA = 1'b0;
            15'b11001101_1001_001: DATA = 1'b0;
            15'b11001101_1001_010: DATA = 1'b0;
            15'b11001101_1001_011: DATA = 1'b0;
            15'b11001101_1001_100: DATA = 1'b1;
            15'b11001101_1001_101: DATA = 1'b1;
            15'b11001101_1001_110: DATA = 1'b0;
            15'b11001101_1001_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 3 Row 10
            15'b11001101_1010_000: DATA = 1'b0;
            15'b11001101_1010_001: DATA = 1'b0;
            15'b11001101_1010_010: DATA = 1'b0;
            15'b11001101_1010_011: DATA = 1'b1;
            15'b11001101_1010_100: DATA = 1'b1;
            15'b11001101_1010_101: DATA = 1'b0;
            15'b11001101_1010_110: DATA = 1'b0;
            15'b11001101_1010_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 3 Row 11
            15'b11001101_1011_000: DATA = 1'b0;
            15'b11001101_1011_001: DATA = 1'b0;
            15'b11001101_1011_010: DATA = 1'b1;
            15'b11001101_1011_011: DATA = 1'b1;
            15'b11001101_1011_100: DATA = 1'b0;
            15'b11001101_1011_101: DATA = 1'b0;
            15'b11001101_1011_110: DATA = 1'b0;
            15'b11001101_1011_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 3 Row 12
            15'b11001101_1100_000: DATA = 1'b1;
            15'b11001101_1100_001: DATA = 1'b1;
            15'b11001101_1100_010: DATA = 1'b1;
            15'b11001101_1100_011: DATA = 1'b0;
            15'b11001101_1100_100: DATA = 1'b0;
            15'b11001101_1100_101: DATA = 1'b0;
            15'b11001101_1100_110: DATA = 1'b0;
            15'b11001101_1100_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 3 Row 13
            15'b11001101_1101_000: DATA = 1'b1;
            15'b11001101_1101_001: DATA = 1'b0;
            15'b11001101_1101_010: DATA = 1'b0;
            15'b11001101_1101_011: DATA = 1'b0;
            15'b11001101_1101_100: DATA = 1'b0;
            15'b11001101_1101_101: DATA = 1'b0;
            15'b11001101_1101_110: DATA = 1'b0;
            15'b11001101_1101_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 3 Row 14
            15'b11001101_1110_000: DATA = 1'b0;
            15'b11001101_1110_001: DATA = 1'b0;
            15'b11001101_1110_010: DATA = 1'b0;
            15'b11001101_1110_011: DATA = 1'b0;
            15'b11001101_1110_100: DATA = 1'b0;
            15'b11001101_1110_101: DATA = 1'b0;
            15'b11001101_1110_110: DATA = 1'b0;
            15'b11001101_1110_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 3 Row 15
            15'b11001101_1111_000: DATA = 1'b0;
            15'b11001101_1111_001: DATA = 1'b0;
            15'b11001101_1111_010: DATA = 1'b0;
            15'b11001101_1111_011: DATA = 1'b0;
            15'b11001101_1111_100: DATA = 1'b0;
            15'b11001101_1111_101: DATA = 1'b0;
            15'b11001101_1111_110: DATA = 1'b0;
            15'b11001101_1111_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 4 Row 0
            15'b11001110_0000_000: DATA = 1'b0;
            15'b11001110_0000_001: DATA = 1'b0;
            15'b11001110_0000_010: DATA = 1'b0;
            15'b11001110_0000_011: DATA = 1'b0;
            15'b11001110_0000_100: DATA = 1'b0;
            15'b11001110_0000_101: DATA = 1'b0;
            15'b11001110_0000_110: DATA = 1'b0;
            15'b11001110_0000_111: DATA = 1'b1;
            //SAWTOOTH- ROW 0 COL 4 Row 1
            15'b11001110_0001_000: DATA = 1'b0;
            15'b11001110_0001_001: DATA = 1'b0;
            15'b11001110_0001_010: DATA = 1'b0;
            15'b11001110_0001_011: DATA = 1'b0;
            15'b11001110_0001_100: DATA = 1'b0;
            15'b11001110_0001_101: DATA = 1'b0;
            15'b11001110_0001_110: DATA = 1'b1;
            15'b11001110_0001_111: DATA = 1'b1;
            //SAWTOOTH- ROW 0 COL 4 Row 2
            15'b11001110_0010_000: DATA = 1'b0;
            15'b11001110_0010_001: DATA = 1'b0;
            15'b11001110_0010_010: DATA = 1'b0;
            15'b11001110_0010_011: DATA = 1'b0;
            15'b11001110_0010_100: DATA = 1'b0;
            15'b11001110_0010_101: DATA = 1'b1;
            15'b11001110_0010_110: DATA = 1'b1;
            15'b11001110_0010_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 4 Row 3
            15'b11001110_0011_000: DATA = 1'b0;
            15'b11001110_0011_001: DATA = 1'b0;
            15'b11001110_0011_010: DATA = 1'b0;
            15'b11001110_0011_011: DATA = 1'b0;
            15'b11001110_0011_100: DATA = 1'b1;
            15'b11001110_0011_101: DATA = 1'b1;
            15'b11001110_0011_110: DATA = 1'b0;
            15'b11001110_0011_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 4 Row 4
            15'b11001110_0100_000: DATA = 1'b0;
            15'b11001110_0100_001: DATA = 1'b0;
            15'b11001110_0100_010: DATA = 1'b1;
            15'b11001110_0100_011: DATA = 1'b1;
            15'b11001110_0100_100: DATA = 1'b1;
            15'b11001110_0100_101: DATA = 1'b0;
            15'b11001110_0100_110: DATA = 1'b0;
            15'b11001110_0100_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 4 Row 5
            15'b11001110_0101_000: DATA = 1'b0;
            15'b11001110_0101_001: DATA = 1'b1;
            15'b11001110_0101_010: DATA = 1'b1;
            15'b11001110_0101_011: DATA = 1'b0;
            15'b11001110_0101_100: DATA = 1'b0;
            15'b11001110_0101_101: DATA = 1'b0;
            15'b11001110_0101_110: DATA = 1'b0;
            15'b11001110_0101_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 4 Row 6
            15'b11001110_0110_000: DATA = 1'b1;
            15'b11001110_0110_001: DATA = 1'b1;
            15'b11001110_0110_010: DATA = 1'b0;
            15'b11001110_0110_011: DATA = 1'b0;
            15'b11001110_0110_100: DATA = 1'b0;
            15'b11001110_0110_101: DATA = 1'b0;
            15'b11001110_0110_110: DATA = 1'b0;
            15'b11001110_0110_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 4 Row 7
            15'b11001110_0111_000: DATA = 1'b1;
            15'b11001110_0111_001: DATA = 1'b0;
            15'b11001110_0111_010: DATA = 1'b0;
            15'b11001110_0111_011: DATA = 1'b0;
            15'b11001110_0111_100: DATA = 1'b0;
            15'b11001110_0111_101: DATA = 1'b0;
            15'b11001110_0111_110: DATA = 1'b0;
            15'b11001110_0111_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 4 Row 8
            15'b11001110_1000_000: DATA = 1'b0;
            15'b11001110_1000_001: DATA = 1'b0;
            15'b11001110_1000_010: DATA = 1'b0;
            15'b11001110_1000_011: DATA = 1'b0;
            15'b11001110_1000_100: DATA = 1'b0;
            15'b11001110_1000_101: DATA = 1'b0;
            15'b11001110_1000_110: DATA = 1'b0;
            15'b11001110_1000_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 4 Row 9
            15'b11001110_1001_000: DATA = 1'b0;
            15'b11001110_1001_001: DATA = 1'b0;
            15'b11001110_1001_010: DATA = 1'b0;
            15'b11001110_1001_011: DATA = 1'b0;
            15'b11001110_1001_100: DATA = 1'b0;
            15'b11001110_1001_101: DATA = 1'b0;
            15'b11001110_1001_110: DATA = 1'b0;
            15'b11001110_1001_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 4 Row 10
            15'b11001110_1010_000: DATA = 1'b0;
            15'b11001110_1010_001: DATA = 1'b0;
            15'b11001110_1010_010: DATA = 1'b0;
            15'b11001110_1010_011: DATA = 1'b0;
            15'b11001110_1010_100: DATA = 1'b0;
            15'b11001110_1010_101: DATA = 1'b0;
            15'b11001110_1010_110: DATA = 1'b0;
            15'b11001110_1010_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 4 Row 11
            15'b11001110_1011_000: DATA = 1'b0;
            15'b11001110_1011_001: DATA = 1'b0;
            15'b11001110_1011_010: DATA = 1'b0;
            15'b11001110_1011_011: DATA = 1'b0;
            15'b11001110_1011_100: DATA = 1'b0;
            15'b11001110_1011_101: DATA = 1'b0;
            15'b11001110_1011_110: DATA = 1'b0;
            15'b11001110_1011_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 4 Row 12
            15'b11001110_1100_000: DATA = 1'b0;
            15'b11001110_1100_001: DATA = 1'b0;
            15'b11001110_1100_010: DATA = 1'b0;
            15'b11001110_1100_011: DATA = 1'b0;
            15'b11001110_1100_100: DATA = 1'b0;
            15'b11001110_1100_101: DATA = 1'b0;
            15'b11001110_1100_110: DATA = 1'b0;
            15'b11001110_1100_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 4 Row 13
            15'b11001110_1101_000: DATA = 1'b0;
            15'b11001110_1101_001: DATA = 1'b0;
            15'b11001110_1101_010: DATA = 1'b0;
            15'b11001110_1101_011: DATA = 1'b0;
            15'b11001110_1101_100: DATA = 1'b0;
            15'b11001110_1101_101: DATA = 1'b0;
            15'b11001110_1101_110: DATA = 1'b0;
            15'b11001110_1101_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 4 Row 14
            15'b11001110_1110_000: DATA = 1'b0;
            15'b11001110_1110_001: DATA = 1'b0;
            15'b11001110_1110_010: DATA = 1'b0;
            15'b11001110_1110_011: DATA = 1'b0;
            15'b11001110_1110_100: DATA = 1'b0;
            15'b11001110_1110_101: DATA = 1'b0;
            15'b11001110_1110_110: DATA = 1'b0;
            15'b11001110_1110_111: DATA = 1'b0;
            //SAWTOOTH- ROW 0 COL 4 Row 15
            15'b11001110_1111_000: DATA = 1'b0;
            15'b11001110_1111_001: DATA = 1'b0;
            15'b11001110_1111_010: DATA = 1'b0;
            15'b11001110_1111_011: DATA = 1'b0;
            15'b11001110_1111_100: DATA = 1'b0;
            15'b11001110_1111_101: DATA = 1'b0;
            15'b11001110_1111_110: DATA = 1'b0;
            15'b11001110_1111_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 0 Row 0
            15'b11001111_0000_000: DATA = 1'b1;
            15'b11001111_0000_001: DATA = 1'b0;
            15'b11001111_0000_010: DATA = 1'b0;
            15'b11001111_0000_011: DATA = 1'b0;
            15'b11001111_0000_100: DATA = 1'b0;
            15'b11001111_0000_101: DATA = 1'b0;
            15'b11001111_0000_110: DATA = 1'b0;
            15'b11001111_0000_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 0 Row 1
            15'b11001111_0001_000: DATA = 1'b1;
            15'b11001111_0001_001: DATA = 1'b0;
            15'b11001111_0001_010: DATA = 1'b0;
            15'b11001111_0001_011: DATA = 1'b0;
            15'b11001111_0001_100: DATA = 1'b0;
            15'b11001111_0001_101: DATA = 1'b0;
            15'b11001111_0001_110: DATA = 1'b0;
            15'b11001111_0001_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 0 Row 2
            15'b11001111_0010_000: DATA = 1'b1;
            15'b11001111_0010_001: DATA = 1'b0;
            15'b11001111_0010_010: DATA = 1'b0;
            15'b11001111_0010_011: DATA = 1'b0;
            15'b11001111_0010_100: DATA = 1'b0;
            15'b11001111_0010_101: DATA = 1'b0;
            15'b11001111_0010_110: DATA = 1'b0;
            15'b11001111_0010_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 0 Row 3
            15'b11001111_0011_000: DATA = 1'b1;
            15'b11001111_0011_001: DATA = 1'b0;
            15'b11001111_0011_010: DATA = 1'b0;
            15'b11001111_0011_011: DATA = 1'b0;
            15'b11001111_0011_100: DATA = 1'b0;
            15'b11001111_0011_101: DATA = 1'b0;
            15'b11001111_0011_110: DATA = 1'b0;
            15'b11001111_0011_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 0 Row 4
            15'b11001111_0100_000: DATA = 1'b1;
            15'b11001111_0100_001: DATA = 1'b0;
            15'b11001111_0100_010: DATA = 1'b0;
            15'b11001111_0100_011: DATA = 1'b0;
            15'b11001111_0100_100: DATA = 1'b0;
            15'b11001111_0100_101: DATA = 1'b0;
            15'b11001111_0100_110: DATA = 1'b0;
            15'b11001111_0100_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 0 Row 5
            15'b11001111_0101_000: DATA = 1'b1;
            15'b11001111_0101_001: DATA = 1'b0;
            15'b11001111_0101_010: DATA = 1'b0;
            15'b11001111_0101_011: DATA = 1'b0;
            15'b11001111_0101_100: DATA = 1'b0;
            15'b11001111_0101_101: DATA = 1'b0;
            15'b11001111_0101_110: DATA = 1'b0;
            15'b11001111_0101_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 0 Row 6
            15'b11001111_0110_000: DATA = 1'b1;
            15'b11001111_0110_001: DATA = 1'b0;
            15'b11001111_0110_010: DATA = 1'b0;
            15'b11001111_0110_011: DATA = 1'b0;
            15'b11001111_0110_100: DATA = 1'b0;
            15'b11001111_0110_101: DATA = 1'b0;
            15'b11001111_0110_110: DATA = 1'b0;
            15'b11001111_0110_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 0 Row 7
            15'b11001111_0111_000: DATA = 1'b1;
            15'b11001111_0111_001: DATA = 1'b0;
            15'b11001111_0111_010: DATA = 1'b0;
            15'b11001111_0111_011: DATA = 1'b0;
            15'b11001111_0111_100: DATA = 1'b0;
            15'b11001111_0111_101: DATA = 1'b0;
            15'b11001111_0111_110: DATA = 1'b0;
            15'b11001111_0111_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 0 Row 8
            15'b11001111_1000_000: DATA = 1'b1;
            15'b11001111_1000_001: DATA = 1'b0;
            15'b11001111_1000_010: DATA = 1'b0;
            15'b11001111_1000_011: DATA = 1'b0;
            15'b11001111_1000_100: DATA = 1'b0;
            15'b11001111_1000_101: DATA = 1'b0;
            15'b11001111_1000_110: DATA = 1'b0;
            15'b11001111_1000_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 0 Row 9
            15'b11001111_1001_000: DATA = 1'b1;
            15'b11001111_1001_001: DATA = 1'b0;
            15'b11001111_1001_010: DATA = 1'b0;
            15'b11001111_1001_011: DATA = 1'b0;
            15'b11001111_1001_100: DATA = 1'b0;
            15'b11001111_1001_101: DATA = 1'b0;
            15'b11001111_1001_110: DATA = 1'b0;
            15'b11001111_1001_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 0 Row 10
            15'b11001111_1010_000: DATA = 1'b1;
            15'b11001111_1010_001: DATA = 1'b0;
            15'b11001111_1010_010: DATA = 1'b0;
            15'b11001111_1010_011: DATA = 1'b0;
            15'b11001111_1010_100: DATA = 1'b0;
            15'b11001111_1010_101: DATA = 1'b0;
            15'b11001111_1010_110: DATA = 1'b0;
            15'b11001111_1010_111: DATA = 1'b1;
            //SAWTOOTH- ROW 1 COL 0 Row 11
            15'b11001111_1011_000: DATA = 1'b1;
            15'b11001111_1011_001: DATA = 1'b0;
            15'b11001111_1011_010: DATA = 1'b0;
            15'b11001111_1011_011: DATA = 1'b0;
            15'b11001111_1011_100: DATA = 1'b0;
            15'b11001111_1011_101: DATA = 1'b0;
            15'b11001111_1011_110: DATA = 1'b1;
            15'b11001111_1011_111: DATA = 1'b1;
            //SAWTOOTH- ROW 1 COL 0 Row 12
            15'b11001111_1100_000: DATA = 1'b1;
            15'b11001111_1100_001: DATA = 1'b0;
            15'b11001111_1100_010: DATA = 1'b0;
            15'b11001111_1100_011: DATA = 1'b0;
            15'b11001111_1100_100: DATA = 1'b1;
            15'b11001111_1100_101: DATA = 1'b1;
            15'b11001111_1100_110: DATA = 1'b1;
            15'b11001111_1100_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 0 Row 13
            15'b11001111_1101_000: DATA = 1'b1;
            15'b11001111_1101_001: DATA = 1'b0;
            15'b11001111_1101_010: DATA = 1'b0;
            15'b11001111_1101_011: DATA = 1'b1;
            15'b11001111_1101_100: DATA = 1'b1;
            15'b11001111_1101_101: DATA = 1'b0;
            15'b11001111_1101_110: DATA = 1'b0;
            15'b11001111_1101_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 0 Row 14
            15'b11001111_1110_000: DATA = 1'b1;
            15'b11001111_1110_001: DATA = 1'b0;
            15'b11001111_1110_010: DATA = 1'b1;
            15'b11001111_1110_011: DATA = 1'b1;
            15'b11001111_1110_100: DATA = 1'b0;
            15'b11001111_1110_101: DATA = 1'b0;
            15'b11001111_1110_110: DATA = 1'b0;
            15'b11001111_1110_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 0 Row 15
            15'b11001111_1111_000: DATA = 1'b1;
            15'b11001111_1111_001: DATA = 1'b1;
            15'b11001111_1111_010: DATA = 1'b0;
            15'b11001111_1111_011: DATA = 1'b0;
            15'b11001111_1111_100: DATA = 1'b0;
            15'b11001111_1111_101: DATA = 1'b0;
            15'b11001111_1111_110: DATA = 1'b0;
            15'b11001111_1111_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 1 Row 0
            15'b11010000_0000_000: DATA = 1'b0;
            15'b11010000_0000_001: DATA = 1'b0;
            15'b11010000_0000_010: DATA = 1'b0;
            15'b11010000_0000_011: DATA = 1'b0;
            15'b11010000_0000_100: DATA = 1'b0;
            15'b11010000_0000_101: DATA = 1'b0;
            15'b11010000_0000_110: DATA = 1'b0;
            15'b11010000_0000_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 1 Row 1
            15'b11010000_0001_000: DATA = 1'b0;
            15'b11010000_0001_001: DATA = 1'b0;
            15'b11010000_0001_010: DATA = 1'b0;
            15'b11010000_0001_011: DATA = 1'b0;
            15'b11010000_0001_100: DATA = 1'b0;
            15'b11010000_0001_101: DATA = 1'b0;
            15'b11010000_0001_110: DATA = 1'b0;
            15'b11010000_0001_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 1 Row 2
            15'b11010000_0010_000: DATA = 1'b0;
            15'b11010000_0010_001: DATA = 1'b0;
            15'b11010000_0010_010: DATA = 1'b0;
            15'b11010000_0010_011: DATA = 1'b0;
            15'b11010000_0010_100: DATA = 1'b0;
            15'b11010000_0010_101: DATA = 1'b0;
            15'b11010000_0010_110: DATA = 1'b0;
            15'b11010000_0010_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 1 Row 3
            15'b11010000_0011_000: DATA = 1'b0;
            15'b11010000_0011_001: DATA = 1'b0;
            15'b11010000_0011_010: DATA = 1'b0;
            15'b11010000_0011_011: DATA = 1'b0;
            15'b11010000_0011_100: DATA = 1'b0;
            15'b11010000_0011_101: DATA = 1'b0;
            15'b11010000_0011_110: DATA = 1'b0;
            15'b11010000_0011_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 1 Row 4
            15'b11010000_0100_000: DATA = 1'b0;
            15'b11010000_0100_001: DATA = 1'b0;
            15'b11010000_0100_010: DATA = 1'b0;
            15'b11010000_0100_011: DATA = 1'b0;
            15'b11010000_0100_100: DATA = 1'b0;
            15'b11010000_0100_101: DATA = 1'b0;
            15'b11010000_0100_110: DATA = 1'b1;
            15'b11010000_0100_111: DATA = 1'b1;
            //SAWTOOTH- ROW 1 COL 1 Row 5
            15'b11010000_0101_000: DATA = 1'b0;
            15'b11010000_0101_001: DATA = 1'b0;
            15'b11010000_0101_010: DATA = 1'b0;
            15'b11010000_0101_011: DATA = 1'b0;
            15'b11010000_0101_100: DATA = 1'b0;
            15'b11010000_0101_101: DATA = 1'b1;
            15'b11010000_0101_110: DATA = 1'b1;
            15'b11010000_0101_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 1 Row 6
            15'b11010000_0110_000: DATA = 1'b0;
            15'b11010000_0110_001: DATA = 1'b0;
            15'b11010000_0110_010: DATA = 1'b0;
            15'b11010000_0110_011: DATA = 1'b0;
            15'b11010000_0110_100: DATA = 1'b1;
            15'b11010000_0110_101: DATA = 1'b1;
            15'b11010000_0110_110: DATA = 1'b0;
            15'b11010000_0110_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 1 Row 7
            15'b11010000_0111_000: DATA = 1'b0;
            15'b11010000_0111_001: DATA = 1'b0;
            15'b11010000_0111_010: DATA = 1'b0;
            15'b11010000_0111_011: DATA = 1'b1;
            15'b11010000_0111_100: DATA = 1'b1;
            15'b11010000_0111_101: DATA = 1'b0;
            15'b11010000_0111_110: DATA = 1'b0;
            15'b11010000_0111_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 1 Row 8
            15'b11010000_1000_000: DATA = 1'b0;
            15'b11010000_1000_001: DATA = 1'b1;
            15'b11010000_1000_010: DATA = 1'b1;
            15'b11010000_1000_011: DATA = 1'b1;
            15'b11010000_1000_100: DATA = 1'b0;
            15'b11010000_1000_101: DATA = 1'b0;
            15'b11010000_1000_110: DATA = 1'b0;
            15'b11010000_1000_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 1 Row 9
            15'b11010000_1001_000: DATA = 1'b1;
            15'b11010000_1001_001: DATA = 1'b1;
            15'b11010000_1001_010: DATA = 1'b0;
            15'b11010000_1001_011: DATA = 1'b0;
            15'b11010000_1001_100: DATA = 1'b0;
            15'b11010000_1001_101: DATA = 1'b0;
            15'b11010000_1001_110: DATA = 1'b0;
            15'b11010000_1001_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 1 Row 10
            15'b11010000_1010_000: DATA = 1'b1;
            15'b11010000_1010_001: DATA = 1'b0;
            15'b11010000_1010_010: DATA = 1'b0;
            15'b11010000_1010_011: DATA = 1'b0;
            15'b11010000_1010_100: DATA = 1'b0;
            15'b11010000_1010_101: DATA = 1'b0;
            15'b11010000_1010_110: DATA = 1'b0;
            15'b11010000_1010_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 1 Row 11
            15'b11010000_1011_000: DATA = 1'b0;
            15'b11010000_1011_001: DATA = 1'b0;
            15'b11010000_1011_010: DATA = 1'b0;
            15'b11010000_1011_011: DATA = 1'b0;
            15'b11010000_1011_100: DATA = 1'b0;
            15'b11010000_1011_101: DATA = 1'b0;
            15'b11010000_1011_110: DATA = 1'b0;
            15'b11010000_1011_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 1 Row 12
            15'b11010000_1100_000: DATA = 1'b0;
            15'b11010000_1100_001: DATA = 1'b0;
            15'b11010000_1100_010: DATA = 1'b0;
            15'b11010000_1100_011: DATA = 1'b0;
            15'b11010000_1100_100: DATA = 1'b0;
            15'b11010000_1100_101: DATA = 1'b0;
            15'b11010000_1100_110: DATA = 1'b0;
            15'b11010000_1100_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 1 Row 13
            15'b11010000_1101_000: DATA = 1'b0;
            15'b11010000_1101_001: DATA = 1'b0;
            15'b11010000_1101_010: DATA = 1'b0;
            15'b11010000_1101_011: DATA = 1'b0;
            15'b11010000_1101_100: DATA = 1'b0;
            15'b11010000_1101_101: DATA = 1'b0;
            15'b11010000_1101_110: DATA = 1'b0;
            15'b11010000_1101_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 1 Row 14
            15'b11010000_1110_000: DATA = 1'b0;
            15'b11010000_1110_001: DATA = 1'b0;
            15'b11010000_1110_010: DATA = 1'b0;
            15'b11010000_1110_011: DATA = 1'b0;
            15'b11010000_1110_100: DATA = 1'b0;
            15'b11010000_1110_101: DATA = 1'b0;
            15'b11010000_1110_110: DATA = 1'b0;
            15'b11010000_1110_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 1 Row 15
            15'b11010000_1111_000: DATA = 1'b0;
            15'b11010000_1111_001: DATA = 1'b0;
            15'b11010000_1111_010: DATA = 1'b0;
            15'b11010000_1111_011: DATA = 1'b0;
            15'b11010000_1111_100: DATA = 1'b0;
            15'b11010000_1111_101: DATA = 1'b0;
            15'b11010000_1111_110: DATA = 1'b0;
            15'b11010000_1111_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 2 Row 0
            15'b11010001_0000_000: DATA = 1'b0;
            15'b11010001_0000_001: DATA = 1'b0;
            15'b11010001_0000_010: DATA = 1'b0;
            15'b11010001_0000_011: DATA = 1'b1;
            15'b11010001_0000_100: DATA = 1'b1;
            15'b11010001_0000_101: DATA = 1'b1;
            15'b11010001_0000_110: DATA = 1'b0;
            15'b11010001_0000_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 2 Row 1
            15'b11010001_0001_000: DATA = 1'b0;
            15'b11010001_0001_001: DATA = 1'b0;
            15'b11010001_0001_010: DATA = 1'b1;
            15'b11010001_0001_011: DATA = 1'b1;
            15'b11010001_0001_100: DATA = 1'b0;
            15'b11010001_0001_101: DATA = 1'b0;
            15'b11010001_0001_110: DATA = 1'b0;
            15'b11010001_0001_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 2 Row 2
            15'b11010001_0010_000: DATA = 1'b0;
            15'b11010001_0010_001: DATA = 1'b1;
            15'b11010001_0010_010: DATA = 1'b1;
            15'b11010001_0010_011: DATA = 1'b0;
            15'b11010001_0010_100: DATA = 1'b0;
            15'b11010001_0010_101: DATA = 1'b0;
            15'b11010001_0010_110: DATA = 1'b0;
            15'b11010001_0010_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 2 Row 3
            15'b11010001_0011_000: DATA = 1'b1;
            15'b11010001_0011_001: DATA = 1'b1;
            15'b11010001_0011_010: DATA = 1'b0;
            15'b11010001_0011_011: DATA = 1'b0;
            15'b11010001_0011_100: DATA = 1'b0;
            15'b11010001_0011_101: DATA = 1'b0;
            15'b11010001_0011_110: DATA = 1'b0;
            15'b11010001_0011_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 2 Row 4
            15'b11010001_0100_000: DATA = 1'b1;
            15'b11010001_0100_001: DATA = 1'b0;
            15'b11010001_0100_010: DATA = 1'b0;
            15'b11010001_0100_011: DATA = 1'b0;
            15'b11010001_0100_100: DATA = 1'b0;
            15'b11010001_0100_101: DATA = 1'b0;
            15'b11010001_0100_110: DATA = 1'b0;
            15'b11010001_0100_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 2 Row 5
            15'b11010001_0101_000: DATA = 1'b0;
            15'b11010001_0101_001: DATA = 1'b0;
            15'b11010001_0101_010: DATA = 1'b0;
            15'b11010001_0101_011: DATA = 1'b0;
            15'b11010001_0101_100: DATA = 1'b0;
            15'b11010001_0101_101: DATA = 1'b0;
            15'b11010001_0101_110: DATA = 1'b0;
            15'b11010001_0101_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 2 Row 6
            15'b11010001_0110_000: DATA = 1'b0;
            15'b11010001_0110_001: DATA = 1'b0;
            15'b11010001_0110_010: DATA = 1'b0;
            15'b11010001_0110_011: DATA = 1'b0;
            15'b11010001_0110_100: DATA = 1'b0;
            15'b11010001_0110_101: DATA = 1'b0;
            15'b11010001_0110_110: DATA = 1'b0;
            15'b11010001_0110_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 2 Row 7
            15'b11010001_0111_000: DATA = 1'b0;
            15'b11010001_0111_001: DATA = 1'b0;
            15'b11010001_0111_010: DATA = 1'b0;
            15'b11010001_0111_011: DATA = 1'b0;
            15'b11010001_0111_100: DATA = 1'b0;
            15'b11010001_0111_101: DATA = 1'b0;
            15'b11010001_0111_110: DATA = 1'b0;
            15'b11010001_0111_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 2 Row 8
            15'b11010001_1000_000: DATA = 1'b0;
            15'b11010001_1000_001: DATA = 1'b0;
            15'b11010001_1000_010: DATA = 1'b0;
            15'b11010001_1000_011: DATA = 1'b0;
            15'b11010001_1000_100: DATA = 1'b0;
            15'b11010001_1000_101: DATA = 1'b0;
            15'b11010001_1000_110: DATA = 1'b0;
            15'b11010001_1000_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 2 Row 9
            15'b11010001_1001_000: DATA = 1'b0;
            15'b11010001_1001_001: DATA = 1'b0;
            15'b11010001_1001_010: DATA = 1'b0;
            15'b11010001_1001_011: DATA = 1'b0;
            15'b11010001_1001_100: DATA = 1'b0;
            15'b11010001_1001_101: DATA = 1'b0;
            15'b11010001_1001_110: DATA = 1'b0;
            15'b11010001_1001_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 2 Row 10
            15'b11010001_1010_000: DATA = 1'b0;
            15'b11010001_1010_001: DATA = 1'b0;
            15'b11010001_1010_010: DATA = 1'b0;
            15'b11010001_1010_011: DATA = 1'b0;
            15'b11010001_1010_100: DATA = 1'b0;
            15'b11010001_1010_101: DATA = 1'b0;
            15'b11010001_1010_110: DATA = 1'b0;
            15'b11010001_1010_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 2 Row 11
            15'b11010001_1011_000: DATA = 1'b0;
            15'b11010001_1011_001: DATA = 1'b0;
            15'b11010001_1011_010: DATA = 1'b0;
            15'b11010001_1011_011: DATA = 1'b0;
            15'b11010001_1011_100: DATA = 1'b0;
            15'b11010001_1011_101: DATA = 1'b0;
            15'b11010001_1011_110: DATA = 1'b0;
            15'b11010001_1011_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 2 Row 12
            15'b11010001_1100_000: DATA = 1'b0;
            15'b11010001_1100_001: DATA = 1'b0;
            15'b11010001_1100_010: DATA = 1'b0;
            15'b11010001_1100_011: DATA = 1'b0;
            15'b11010001_1100_100: DATA = 1'b0;
            15'b11010001_1100_101: DATA = 1'b0;
            15'b11010001_1100_110: DATA = 1'b0;
            15'b11010001_1100_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 2 Row 13
            15'b11010001_1101_000: DATA = 1'b0;
            15'b11010001_1101_001: DATA = 1'b0;
            15'b11010001_1101_010: DATA = 1'b0;
            15'b11010001_1101_011: DATA = 1'b0;
            15'b11010001_1101_100: DATA = 1'b0;
            15'b11010001_1101_101: DATA = 1'b0;
            15'b11010001_1101_110: DATA = 1'b0;
            15'b11010001_1101_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 2 Row 14
            15'b11010001_1110_000: DATA = 1'b0;
            15'b11010001_1110_001: DATA = 1'b0;
            15'b11010001_1110_010: DATA = 1'b0;
            15'b11010001_1110_011: DATA = 1'b0;
            15'b11010001_1110_100: DATA = 1'b0;
            15'b11010001_1110_101: DATA = 1'b0;
            15'b11010001_1110_110: DATA = 1'b0;
            15'b11010001_1110_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 2 Row 15
            15'b11010001_1111_000: DATA = 1'b0;
            15'b11010001_1111_001: DATA = 1'b0;
            15'b11010001_1111_010: DATA = 1'b0;
            15'b11010001_1111_011: DATA = 1'b0;
            15'b11010001_1111_100: DATA = 1'b0;
            15'b11010001_1111_101: DATA = 1'b0;
            15'b11010001_1111_110: DATA = 1'b0;
            15'b11010001_1111_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 3 Row 0
            15'b11010010_0000_000: DATA = 1'b0;
            15'b11010010_0000_001: DATA = 1'b0;
            15'b11010010_0000_010: DATA = 1'b0;
            15'b11010010_0000_011: DATA = 1'b0;
            15'b11010010_0000_100: DATA = 1'b0;
            15'b11010010_0000_101: DATA = 1'b0;
            15'b11010010_0000_110: DATA = 1'b0;
            15'b11010010_0000_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 3 Row 1
            15'b11010010_0001_000: DATA = 1'b0;
            15'b11010010_0001_001: DATA = 1'b0;
            15'b11010010_0001_010: DATA = 1'b0;
            15'b11010010_0001_011: DATA = 1'b0;
            15'b11010010_0001_100: DATA = 1'b0;
            15'b11010010_0001_101: DATA = 1'b0;
            15'b11010010_0001_110: DATA = 1'b0;
            15'b11010010_0001_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 3 Row 2
            15'b11010010_0010_000: DATA = 1'b0;
            15'b11010010_0010_001: DATA = 1'b0;
            15'b11010010_0010_010: DATA = 1'b0;
            15'b11010010_0010_011: DATA = 1'b0;
            15'b11010010_0010_100: DATA = 1'b0;
            15'b11010010_0010_101: DATA = 1'b0;
            15'b11010010_0010_110: DATA = 1'b0;
            15'b11010010_0010_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 3 Row 3
            15'b11010010_0011_000: DATA = 1'b0;
            15'b11010010_0011_001: DATA = 1'b0;
            15'b11010010_0011_010: DATA = 1'b0;
            15'b11010010_0011_011: DATA = 1'b0;
            15'b11010010_0011_100: DATA = 1'b0;
            15'b11010010_0011_101: DATA = 1'b0;
            15'b11010010_0011_110: DATA = 1'b0;
            15'b11010010_0011_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 3 Row 4
            15'b11010010_0100_000: DATA = 1'b0;
            15'b11010010_0100_001: DATA = 1'b0;
            15'b11010010_0100_010: DATA = 1'b0;
            15'b11010010_0100_011: DATA = 1'b0;
            15'b11010010_0100_100: DATA = 1'b0;
            15'b11010010_0100_101: DATA = 1'b0;
            15'b11010010_0100_110: DATA = 1'b0;
            15'b11010010_0100_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 3 Row 5
            15'b11010010_0101_000: DATA = 1'b0;
            15'b11010010_0101_001: DATA = 1'b0;
            15'b11010010_0101_010: DATA = 1'b0;
            15'b11010010_0101_011: DATA = 1'b0;
            15'b11010010_0101_100: DATA = 1'b0;
            15'b11010010_0101_101: DATA = 1'b0;
            15'b11010010_0101_110: DATA = 1'b0;
            15'b11010010_0101_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 3 Row 6
            15'b11010010_0110_000: DATA = 1'b0;
            15'b11010010_0110_001: DATA = 1'b0;
            15'b11010010_0110_010: DATA = 1'b0;
            15'b11010010_0110_011: DATA = 1'b0;
            15'b11010010_0110_100: DATA = 1'b0;
            15'b11010010_0110_101: DATA = 1'b0;
            15'b11010010_0110_110: DATA = 1'b0;
            15'b11010010_0110_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 3 Row 7
            15'b11010010_0111_000: DATA = 1'b0;
            15'b11010010_0111_001: DATA = 1'b0;
            15'b11010010_0111_010: DATA = 1'b0;
            15'b11010010_0111_011: DATA = 1'b0;
            15'b11010010_0111_100: DATA = 1'b0;
            15'b11010010_0111_101: DATA = 1'b0;
            15'b11010010_0111_110: DATA = 1'b0;
            15'b11010010_0111_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 3 Row 8
            15'b11010010_1000_000: DATA = 1'b0;
            15'b11010010_1000_001: DATA = 1'b0;
            15'b11010010_1000_010: DATA = 1'b0;
            15'b11010010_1000_011: DATA = 1'b0;
            15'b11010010_1000_100: DATA = 1'b0;
            15'b11010010_1000_101: DATA = 1'b0;
            15'b11010010_1000_110: DATA = 1'b0;
            15'b11010010_1000_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 3 Row 9
            15'b11010010_1001_000: DATA = 1'b0;
            15'b11010010_1001_001: DATA = 1'b0;
            15'b11010010_1001_010: DATA = 1'b0;
            15'b11010010_1001_011: DATA = 1'b0;
            15'b11010010_1001_100: DATA = 1'b0;
            15'b11010010_1001_101: DATA = 1'b0;
            15'b11010010_1001_110: DATA = 1'b0;
            15'b11010010_1001_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 3 Row 10
            15'b11010010_1010_000: DATA = 1'b0;
            15'b11010010_1010_001: DATA = 1'b0;
            15'b11010010_1010_010: DATA = 1'b0;
            15'b11010010_1010_011: DATA = 1'b0;
            15'b11010010_1010_100: DATA = 1'b0;
            15'b11010010_1010_101: DATA = 1'b0;
            15'b11010010_1010_110: DATA = 1'b0;
            15'b11010010_1010_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 3 Row 11
            15'b11010010_1011_000: DATA = 1'b0;
            15'b11010010_1011_001: DATA = 1'b0;
            15'b11010010_1011_010: DATA = 1'b0;
            15'b11010010_1011_011: DATA = 1'b0;
            15'b11010010_1011_100: DATA = 1'b0;
            15'b11010010_1011_101: DATA = 1'b0;
            15'b11010010_1011_110: DATA = 1'b0;
            15'b11010010_1011_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 3 Row 12
            15'b11010010_1100_000: DATA = 1'b0;
            15'b11010010_1100_001: DATA = 1'b0;
            15'b11010010_1100_010: DATA = 1'b0;
            15'b11010010_1100_011: DATA = 1'b0;
            15'b11010010_1100_100: DATA = 1'b0;
            15'b11010010_1100_101: DATA = 1'b0;
            15'b11010010_1100_110: DATA = 1'b0;
            15'b11010010_1100_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 3 Row 13
            15'b11010010_1101_000: DATA = 1'b0;
            15'b11010010_1101_001: DATA = 1'b0;
            15'b11010010_1101_010: DATA = 1'b0;
            15'b11010010_1101_011: DATA = 1'b0;
            15'b11010010_1101_100: DATA = 1'b0;
            15'b11010010_1101_101: DATA = 1'b0;
            15'b11010010_1101_110: DATA = 1'b0;
            15'b11010010_1101_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 3 Row 14
            15'b11010010_1110_000: DATA = 1'b0;
            15'b11010010_1110_001: DATA = 1'b0;
            15'b11010010_1110_010: DATA = 1'b0;
            15'b11010010_1110_011: DATA = 1'b0;
            15'b11010010_1110_100: DATA = 1'b0;
            15'b11010010_1110_101: DATA = 1'b0;
            15'b11010010_1110_110: DATA = 1'b0;
            15'b11010010_1110_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 3 Row 15
            15'b11010010_1111_000: DATA = 1'b0;
            15'b11010010_1111_001: DATA = 1'b0;
            15'b11010010_1111_010: DATA = 1'b0;
            15'b11010010_1111_011: DATA = 1'b0;
            15'b11010010_1111_100: DATA = 1'b0;
            15'b11010010_1111_101: DATA = 1'b0;
            15'b11010010_1111_110: DATA = 1'b0;
            15'b11010010_1111_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 4 Row 0
            15'b11010011_0000_000: DATA = 1'b0;
            15'b11010011_0000_001: DATA = 1'b0;
            15'b11010011_0000_010: DATA = 1'b0;
            15'b11010011_0000_011: DATA = 1'b0;
            15'b11010011_0000_100: DATA = 1'b0;
            15'b11010011_0000_101: DATA = 1'b0;
            15'b11010011_0000_110: DATA = 1'b0;
            15'b11010011_0000_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 4 Row 1
            15'b11010011_0001_000: DATA = 1'b0;
            15'b11010011_0001_001: DATA = 1'b0;
            15'b11010011_0001_010: DATA = 1'b0;
            15'b11010011_0001_011: DATA = 1'b0;
            15'b11010011_0001_100: DATA = 1'b0;
            15'b11010011_0001_101: DATA = 1'b0;
            15'b11010011_0001_110: DATA = 1'b0;
            15'b11010011_0001_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 4 Row 2
            15'b11010011_0010_000: DATA = 1'b0;
            15'b11010011_0010_001: DATA = 1'b0;
            15'b11010011_0010_010: DATA = 1'b0;
            15'b11010011_0010_011: DATA = 1'b0;
            15'b11010011_0010_100: DATA = 1'b0;
            15'b11010011_0010_101: DATA = 1'b0;
            15'b11010011_0010_110: DATA = 1'b0;
            15'b11010011_0010_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 4 Row 3
            15'b11010011_0011_000: DATA = 1'b0;
            15'b11010011_0011_001: DATA = 1'b0;
            15'b11010011_0011_010: DATA = 1'b0;
            15'b11010011_0011_011: DATA = 1'b0;
            15'b11010011_0011_100: DATA = 1'b0;
            15'b11010011_0011_101: DATA = 1'b0;
            15'b11010011_0011_110: DATA = 1'b0;
            15'b11010011_0011_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 4 Row 4
            15'b11010011_0100_000: DATA = 1'b0;
            15'b11010011_0100_001: DATA = 1'b0;
            15'b11010011_0100_010: DATA = 1'b0;
            15'b11010011_0100_011: DATA = 1'b0;
            15'b11010011_0100_100: DATA = 1'b0;
            15'b11010011_0100_101: DATA = 1'b0;
            15'b11010011_0100_110: DATA = 1'b0;
            15'b11010011_0100_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 4 Row 5
            15'b11010011_0101_000: DATA = 1'b0;
            15'b11010011_0101_001: DATA = 1'b0;
            15'b11010011_0101_010: DATA = 1'b0;
            15'b11010011_0101_011: DATA = 1'b0;
            15'b11010011_0101_100: DATA = 1'b0;
            15'b11010011_0101_101: DATA = 1'b0;
            15'b11010011_0101_110: DATA = 1'b0;
            15'b11010011_0101_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 4 Row 6
            15'b11010011_0110_000: DATA = 1'b0;
            15'b11010011_0110_001: DATA = 1'b0;
            15'b11010011_0110_010: DATA = 1'b0;
            15'b11010011_0110_011: DATA = 1'b0;
            15'b11010011_0110_100: DATA = 1'b0;
            15'b11010011_0110_101: DATA = 1'b0;
            15'b11010011_0110_110: DATA = 1'b0;
            15'b11010011_0110_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 4 Row 7
            15'b11010011_0111_000: DATA = 1'b0;
            15'b11010011_0111_001: DATA = 1'b0;
            15'b11010011_0111_010: DATA = 1'b0;
            15'b11010011_0111_011: DATA = 1'b0;
            15'b11010011_0111_100: DATA = 1'b0;
            15'b11010011_0111_101: DATA = 1'b0;
            15'b11010011_0111_110: DATA = 1'b0;
            15'b11010011_0111_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 4 Row 8
            15'b11010011_1000_000: DATA = 1'b0;
            15'b11010011_1000_001: DATA = 1'b0;
            15'b11010011_1000_010: DATA = 1'b0;
            15'b11010011_1000_011: DATA = 1'b0;
            15'b11010011_1000_100: DATA = 1'b0;
            15'b11010011_1000_101: DATA = 1'b0;
            15'b11010011_1000_110: DATA = 1'b0;
            15'b11010011_1000_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 4 Row 9
            15'b11010011_1001_000: DATA = 1'b0;
            15'b11010011_1001_001: DATA = 1'b0;
            15'b11010011_1001_010: DATA = 1'b0;
            15'b11010011_1001_011: DATA = 1'b0;
            15'b11010011_1001_100: DATA = 1'b0;
            15'b11010011_1001_101: DATA = 1'b0;
            15'b11010011_1001_110: DATA = 1'b0;
            15'b11010011_1001_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 4 Row 10
            15'b11010011_1010_000: DATA = 1'b0;
            15'b11010011_1010_001: DATA = 1'b0;
            15'b11010011_1010_010: DATA = 1'b0;
            15'b11010011_1010_011: DATA = 1'b0;
            15'b11010011_1010_100: DATA = 1'b0;
            15'b11010011_1010_101: DATA = 1'b0;
            15'b11010011_1010_110: DATA = 1'b0;
            15'b11010011_1010_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 4 Row 11
            15'b11010011_1011_000: DATA = 1'b0;
            15'b11010011_1011_001: DATA = 1'b0;
            15'b11010011_1011_010: DATA = 1'b0;
            15'b11010011_1011_011: DATA = 1'b0;
            15'b11010011_1011_100: DATA = 1'b0;
            15'b11010011_1011_101: DATA = 1'b0;
            15'b11010011_1011_110: DATA = 1'b0;
            15'b11010011_1011_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 4 Row 12
            15'b11010011_1100_000: DATA = 1'b0;
            15'b11010011_1100_001: DATA = 1'b0;
            15'b11010011_1100_010: DATA = 1'b0;
            15'b11010011_1100_011: DATA = 1'b0;
            15'b11010011_1100_100: DATA = 1'b0;
            15'b11010011_1100_101: DATA = 1'b0;
            15'b11010011_1100_110: DATA = 1'b0;
            15'b11010011_1100_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 4 Row 13
            15'b11010011_1101_000: DATA = 1'b0;
            15'b11010011_1101_001: DATA = 1'b0;
            15'b11010011_1101_010: DATA = 1'b0;
            15'b11010011_1101_011: DATA = 1'b0;
            15'b11010011_1101_100: DATA = 1'b0;
            15'b11010011_1101_101: DATA = 1'b0;
            15'b11010011_1101_110: DATA = 1'b0;
            15'b11010011_1101_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 4 Row 14
            15'b11010011_1110_000: DATA = 1'b0;
            15'b11010011_1110_001: DATA = 1'b0;
            15'b11010011_1110_010: DATA = 1'b0;
            15'b11010011_1110_011: DATA = 1'b0;
            15'b11010011_1110_100: DATA = 1'b0;
            15'b11010011_1110_101: DATA = 1'b0;
            15'b11010011_1110_110: DATA = 1'b0;
            15'b11010011_1110_111: DATA = 1'b0;
            //SAWTOOTH- ROW 1 COL 4 Row 15
            15'b11010011_1111_000: DATA = 1'b0;
            15'b11010011_1111_001: DATA = 1'b0;
            15'b11010011_1111_010: DATA = 1'b0;
            15'b11010011_1111_011: DATA = 1'b0;
            15'b11010011_1111_100: DATA = 1'b0;
            15'b11010011_1111_101: DATA = 1'b0;
            15'b11010011_1111_110: DATA = 1'b0;
            15'b11010011_1111_111: DATA = 1'b0;
            //UPPER LEFT 0 COL 0 Row 0
            15'b11010100_0000_000: DATA = 1'b1;
            15'b11010100_0000_001: DATA = 1'b1;
            15'b11010100_0000_010: DATA = 1'b1;
            15'b11010100_0000_011: DATA = 1'b1;
            15'b11010100_0000_100: DATA = 1'b1;
            15'b11010100_0000_101: DATA = 1'b1;
            15'b11010100_0000_110: DATA = 1'b1;
            15'b11010100_0000_111: DATA = 1'b1;
            //UPPER LEFT 0 COL 0 Row 1
            15'b11010100_0001_000: DATA = 1'b1;
            15'b11010100_0001_001: DATA = 1'b0;
            15'b11010100_0001_010: DATA = 1'b0;
            15'b11010100_0001_011: DATA = 1'b0;
            15'b11010100_0001_100: DATA = 1'b0;
            15'b11010100_0001_101: DATA = 1'b0;
            15'b11010100_0001_110: DATA = 1'b0;
            15'b11010100_0001_111: DATA = 1'b0;
            //UPPER LEFT 0 COL 0 Row 2
            15'b11010100_0010_000: DATA = 1'b1;
            15'b11010100_0010_001: DATA = 1'b0;
            15'b11010100_0010_010: DATA = 1'b0;
            15'b11010100_0010_011: DATA = 1'b0;
            15'b11010100_0010_100: DATA = 1'b0;
            15'b11010100_0010_101: DATA = 1'b0;
            15'b11010100_0010_110: DATA = 1'b0;
            15'b11010100_0010_111: DATA = 1'b0;
            //UPPER LEFT 0 COL 0 Row 3
            15'b11010100_0011_000: DATA = 1'b1;
            15'b11010100_0011_001: DATA = 1'b0;
            15'b11010100_0011_010: DATA = 1'b0;
            15'b11010100_0011_011: DATA = 1'b0;
            15'b11010100_0011_100: DATA = 1'b0;
            15'b11010100_0011_101: DATA = 1'b0;
            15'b11010100_0011_110: DATA = 1'b0;
            15'b11010100_0011_111: DATA = 1'b0;
            //UPPER LEFT 0 COL 0 Row 4
            15'b11010100_0100_000: DATA = 1'b1;
            15'b11010100_0100_001: DATA = 1'b0;
            15'b11010100_0100_010: DATA = 1'b0;
            15'b11010100_0100_011: DATA = 1'b0;
            15'b11010100_0100_100: DATA = 1'b0;
            15'b11010100_0100_101: DATA = 1'b0;
            15'b11010100_0100_110: DATA = 1'b0;
            15'b11010100_0100_111: DATA = 1'b0;
            //UPPER LEFT 0 COL 0 Row 5
            15'b11010100_0101_000: DATA = 1'b1;
            15'b11010100_0101_001: DATA = 1'b0;
            15'b11010100_0101_010: DATA = 1'b0;
            15'b11010100_0101_011: DATA = 1'b0;
            15'b11010100_0101_100: DATA = 1'b0;
            15'b11010100_0101_101: DATA = 1'b0;
            15'b11010100_0101_110: DATA = 1'b0;
            15'b11010100_0101_111: DATA = 1'b0;
            //UPPER LEFT 0 COL 0 Row 6
            15'b11010100_0110_000: DATA = 1'b1;
            15'b11010100_0110_001: DATA = 1'b0;
            15'b11010100_0110_010: DATA = 1'b0;
            15'b11010100_0110_011: DATA = 1'b0;
            15'b11010100_0110_100: DATA = 1'b0;
            15'b11010100_0110_101: DATA = 1'b0;
            15'b11010100_0110_110: DATA = 1'b0;
            15'b11010100_0110_111: DATA = 1'b0;
            //UPPER LEFT 0 COL 0 Row 7
            15'b11010100_0111_000: DATA = 1'b1;
            15'b11010100_0111_001: DATA = 1'b0;
            15'b11010100_0111_010: DATA = 1'b0;
            15'b11010100_0111_011: DATA = 1'b0;
            15'b11010100_0111_100: DATA = 1'b0;
            15'b11010100_0111_101: DATA = 1'b0;
            15'b11010100_0111_110: DATA = 1'b0;
            15'b11010100_0111_111: DATA = 1'b0;
            //UPPER LEFT 0 COL 0 Row 8
            15'b11010100_1000_000: DATA = 1'b1;
            15'b11010100_1000_001: DATA = 1'b0;
            15'b11010100_1000_010: DATA = 1'b0;
            15'b11010100_1000_011: DATA = 1'b0;
            15'b11010100_1000_100: DATA = 1'b0;
            15'b11010100_1000_101: DATA = 1'b0;
            15'b11010100_1000_110: DATA = 1'b0;
            15'b11010100_1000_111: DATA = 1'b0;
            //UPPER LEFT 0 COL 0 Row 9
            15'b11010100_1001_000: DATA = 1'b1;
            15'b11010100_1001_001: DATA = 1'b0;
            15'b11010100_1001_010: DATA = 1'b0;
            15'b11010100_1001_011: DATA = 1'b0;
            15'b11010100_1001_100: DATA = 1'b0;
            15'b11010100_1001_101: DATA = 1'b0;
            15'b11010100_1001_110: DATA = 1'b0;
            15'b11010100_1001_111: DATA = 1'b0;
            //UPPER LEFT 0 COL 0 Row 10
            15'b11010100_1010_000: DATA = 1'b1;
            15'b11010100_1010_001: DATA = 1'b0;
            15'b11010100_1010_010: DATA = 1'b0;
            15'b11010100_1010_011: DATA = 1'b0;
            15'b11010100_1010_100: DATA = 1'b0;
            15'b11010100_1010_101: DATA = 1'b0;
            15'b11010100_1010_110: DATA = 1'b0;
            15'b11010100_1010_111: DATA = 1'b0;
            //UPPER LEFT 0 COL 0 Row 11
            15'b11010100_1011_000: DATA = 1'b1;
            15'b11010100_1011_001: DATA = 1'b0;
            15'b11010100_1011_010: DATA = 1'b0;
            15'b11010100_1011_011: DATA = 1'b0;
            15'b11010100_1011_100: DATA = 1'b0;
            15'b11010100_1011_101: DATA = 1'b0;
            15'b11010100_1011_110: DATA = 1'b0;
            15'b11010100_1011_111: DATA = 1'b0;
            //UPPER LEFT 0 COL 0 Row 12
            15'b11010100_1100_000: DATA = 1'b1;
            15'b11010100_1100_001: DATA = 1'b0;
            15'b11010100_1100_010: DATA = 1'b0;
            15'b11010100_1100_011: DATA = 1'b0;
            15'b11010100_1100_100: DATA = 1'b0;
            15'b11010100_1100_101: DATA = 1'b0;
            15'b11010100_1100_110: DATA = 1'b0;
            15'b11010100_1100_111: DATA = 1'b0;
            //UPPER LEFT 0 COL 0 Row 13
            15'b11010100_1101_000: DATA = 1'b1;
            15'b11010100_1101_001: DATA = 1'b0;
            15'b11010100_1101_010: DATA = 1'b0;
            15'b11010100_1101_011: DATA = 1'b0;
            15'b11010100_1101_100: DATA = 1'b0;
            15'b11010100_1101_101: DATA = 1'b0;
            15'b11010100_1101_110: DATA = 1'b0;
            15'b11010100_1101_111: DATA = 1'b0;
            //UPPER LEFT 0 COL 0 Row 14
            15'b11010100_1110_000: DATA = 1'b1;
            15'b11010100_1110_001: DATA = 1'b0;
            15'b11010100_1110_010: DATA = 1'b0;
            15'b11010100_1110_011: DATA = 1'b0;
            15'b11010100_1110_100: DATA = 1'b0;
            15'b11010100_1110_101: DATA = 1'b0;
            15'b11010100_1110_110: DATA = 1'b0;
            15'b11010100_1110_111: DATA = 1'b0;
            //UPPER LEFT 0 COL 0 Row 15
            15'b11010100_1111_000: DATA = 1'b1;
            15'b11010100_1111_001: DATA = 1'b0;
            15'b11010100_1111_010: DATA = 1'b0;
            15'b11010100_1111_011: DATA = 1'b0;
            15'b11010100_1111_100: DATA = 1'b0;
            15'b11010100_1111_101: DATA = 1'b0;
            15'b11010100_1111_110: DATA = 1'b0;
            15'b11010100_1111_111: DATA = 1'b0;
            //UPPER RIGHT 0 COL 0 Row 0
            15'b11010101_0000_000: DATA = 1'b1;
            15'b11010101_0000_001: DATA = 1'b1;
            15'b11010101_0000_010: DATA = 1'b1;
            15'b11010101_0000_011: DATA = 1'b1;
            15'b11010101_0000_100: DATA = 1'b1;
            15'b11010101_0000_101: DATA = 1'b1;
            15'b11010101_0000_110: DATA = 1'b1;
            15'b11010101_0000_111: DATA = 1'b1;
            //UPPER RIGHT 0 COL 0 Row 1
            15'b11010101_0001_000: DATA = 1'b0;
            15'b11010101_0001_001: DATA = 1'b0;
            15'b11010101_0001_010: DATA = 1'b0;
            15'b11010101_0001_011: DATA = 1'b0;
            15'b11010101_0001_100: DATA = 1'b0;
            15'b11010101_0001_101: DATA = 1'b0;
            15'b11010101_0001_110: DATA = 1'b0;
            15'b11010101_0001_111: DATA = 1'b1;
            //UPPER RIGHT 0 COL 0 Row 2
            15'b11010101_0010_000: DATA = 1'b0;
            15'b11010101_0010_001: DATA = 1'b0;
            15'b11010101_0010_010: DATA = 1'b0;
            15'b11010101_0010_011: DATA = 1'b0;
            15'b11010101_0010_100: DATA = 1'b0;
            15'b11010101_0010_101: DATA = 1'b0;
            15'b11010101_0010_110: DATA = 1'b0;
            15'b11010101_0010_111: DATA = 1'b1;
            //UPPER RIGHT 0 COL 0 Row 3
            15'b11010101_0011_000: DATA = 1'b0;
            15'b11010101_0011_001: DATA = 1'b0;
            15'b11010101_0011_010: DATA = 1'b0;
            15'b11010101_0011_011: DATA = 1'b0;
            15'b11010101_0011_100: DATA = 1'b0;
            15'b11010101_0011_101: DATA = 1'b0;
            15'b11010101_0011_110: DATA = 1'b0;
            15'b11010101_0011_111: DATA = 1'b1;
            //UPPER RIGHT 0 COL 0 Row 4
            15'b11010101_0100_000: DATA = 1'b0;
            15'b11010101_0100_001: DATA = 1'b0;
            15'b11010101_0100_010: DATA = 1'b0;
            15'b11010101_0100_011: DATA = 1'b0;
            15'b11010101_0100_100: DATA = 1'b0;
            15'b11010101_0100_101: DATA = 1'b0;
            15'b11010101_0100_110: DATA = 1'b0;
            15'b11010101_0100_111: DATA = 1'b1;
            //UPPER RIGHT 0 COL 0 Row 5
            15'b11010101_0101_000: DATA = 1'b0;
            15'b11010101_0101_001: DATA = 1'b0;
            15'b11010101_0101_010: DATA = 1'b0;
            15'b11010101_0101_011: DATA = 1'b0;
            15'b11010101_0101_100: DATA = 1'b0;
            15'b11010101_0101_101: DATA = 1'b0;
            15'b11010101_0101_110: DATA = 1'b0;
            15'b11010101_0101_111: DATA = 1'b1;
            //UPPER RIGHT 0 COL 0 Row 6
            15'b11010101_0110_000: DATA = 1'b0;
            15'b11010101_0110_001: DATA = 1'b0;
            15'b11010101_0110_010: DATA = 1'b0;
            15'b11010101_0110_011: DATA = 1'b0;
            15'b11010101_0110_100: DATA = 1'b0;
            15'b11010101_0110_101: DATA = 1'b0;
            15'b11010101_0110_110: DATA = 1'b0;
            15'b11010101_0110_111: DATA = 1'b1;
            //UPPER RIGHT 0 COL 0 Row 7
            15'b11010101_0111_000: DATA = 1'b0;
            15'b11010101_0111_001: DATA = 1'b0;
            15'b11010101_0111_010: DATA = 1'b0;
            15'b11010101_0111_011: DATA = 1'b0;
            15'b11010101_0111_100: DATA = 1'b0;
            15'b11010101_0111_101: DATA = 1'b0;
            15'b11010101_0111_110: DATA = 1'b0;
            15'b11010101_0111_111: DATA = 1'b1;
            //UPPER RIGHT 0 COL 0 Row 8
            15'b11010101_1000_000: DATA = 1'b0;
            15'b11010101_1000_001: DATA = 1'b0;
            15'b11010101_1000_010: DATA = 1'b0;
            15'b11010101_1000_011: DATA = 1'b0;
            15'b11010101_1000_100: DATA = 1'b0;
            15'b11010101_1000_101: DATA = 1'b0;
            15'b11010101_1000_110: DATA = 1'b0;
            15'b11010101_1000_111: DATA = 1'b1;
            //UPPER RIGHT 0 COL 0 Row 9
            15'b11010101_1001_000: DATA = 1'b0;
            15'b11010101_1001_001: DATA = 1'b0;
            15'b11010101_1001_010: DATA = 1'b0;
            15'b11010101_1001_011: DATA = 1'b0;
            15'b11010101_1001_100: DATA = 1'b0;
            15'b11010101_1001_101: DATA = 1'b0;
            15'b11010101_1001_110: DATA = 1'b0;
            15'b11010101_1001_111: DATA = 1'b1;
            //UPPER RIGHT 0 COL 0 Row 10
            15'b11010101_1010_000: DATA = 1'b0;
            15'b11010101_1010_001: DATA = 1'b0;
            15'b11010101_1010_010: DATA = 1'b0;
            15'b11010101_1010_011: DATA = 1'b0;
            15'b11010101_1010_100: DATA = 1'b0;
            15'b11010101_1010_101: DATA = 1'b0;
            15'b11010101_1010_110: DATA = 1'b0;
            15'b11010101_1010_111: DATA = 1'b1;
            //UPPER RIGHT 0 COL 0 Row 11
            15'b11010101_1011_000: DATA = 1'b0;
            15'b11010101_1011_001: DATA = 1'b0;
            15'b11010101_1011_010: DATA = 1'b0;
            15'b11010101_1011_011: DATA = 1'b0;
            15'b11010101_1011_100: DATA = 1'b0;
            15'b11010101_1011_101: DATA = 1'b0;
            15'b11010101_1011_110: DATA = 1'b0;
            15'b11010101_1011_111: DATA = 1'b1;
            //UPPER RIGHT 0 COL 0 Row 12
            15'b11010101_1100_000: DATA = 1'b0;
            15'b11010101_1100_001: DATA = 1'b0;
            15'b11010101_1100_010: DATA = 1'b0;
            15'b11010101_1100_011: DATA = 1'b0;
            15'b11010101_1100_100: DATA = 1'b0;
            15'b11010101_1100_101: DATA = 1'b0;
            15'b11010101_1100_110: DATA = 1'b0;
            15'b11010101_1100_111: DATA = 1'b1;
            //UPPER RIGHT 0 COL 0 Row 13
            15'b11010101_1101_000: DATA = 1'b0;
            15'b11010101_1101_001: DATA = 1'b0;
            15'b11010101_1101_010: DATA = 1'b0;
            15'b11010101_1101_011: DATA = 1'b0;
            15'b11010101_1101_100: DATA = 1'b0;
            15'b11010101_1101_101: DATA = 1'b0;
            15'b11010101_1101_110: DATA = 1'b0;
            15'b11010101_1101_111: DATA = 1'b1;
            //UPPER RIGHT 0 COL 0 Row 14
            15'b11010101_1110_000: DATA = 1'b0;
            15'b11010101_1110_001: DATA = 1'b0;
            15'b11010101_1110_010: DATA = 1'b0;
            15'b11010101_1110_011: DATA = 1'b0;
            15'b11010101_1110_100: DATA = 1'b0;
            15'b11010101_1110_101: DATA = 1'b0;
            15'b11010101_1110_110: DATA = 1'b0;
            15'b11010101_1110_111: DATA = 1'b1;
            //UPPER RIGHT 0 COL 0 Row 15
            15'b11010101_1111_000: DATA = 1'b0;
            15'b11010101_1111_001: DATA = 1'b0;
            15'b11010101_1111_010: DATA = 1'b0;
            15'b11010101_1111_011: DATA = 1'b0;
            15'b11010101_1111_100: DATA = 1'b0;
            15'b11010101_1111_101: DATA = 1'b0;
            15'b11010101_1111_110: DATA = 1'b0;
            15'b11010101_1111_111: DATA = 1'b1;
            //BOTTOM LEFT 0 COL 0 Row 0
            15'b11010110_0000_000: DATA = 1'b1;
            15'b11010110_0000_001: DATA = 1'b0;
            15'b11010110_0000_010: DATA = 1'b0;
            15'b11010110_0000_011: DATA = 1'b0;
            15'b11010110_0000_100: DATA = 1'b0;
            15'b11010110_0000_101: DATA = 1'b0;
            15'b11010110_0000_110: DATA = 1'b0;
            15'b11010110_0000_111: DATA = 1'b0;
            //BOTTOM LEFT 0 COL 0 Row 1
            15'b11010110_0001_000: DATA = 1'b1;
            15'b11010110_0001_001: DATA = 1'b0;
            15'b11010110_0001_010: DATA = 1'b0;
            15'b11010110_0001_011: DATA = 1'b0;
            15'b11010110_0001_100: DATA = 1'b0;
            15'b11010110_0001_101: DATA = 1'b0;
            15'b11010110_0001_110: DATA = 1'b0;
            15'b11010110_0001_111: DATA = 1'b0;
            //BOTTOM LEFT 0 COL 0 Row 2
            15'b11010110_0010_000: DATA = 1'b1;
            15'b11010110_0010_001: DATA = 1'b0;
            15'b11010110_0010_010: DATA = 1'b0;
            15'b11010110_0010_011: DATA = 1'b0;
            15'b11010110_0010_100: DATA = 1'b0;
            15'b11010110_0010_101: DATA = 1'b0;
            15'b11010110_0010_110: DATA = 1'b0;
            15'b11010110_0010_111: DATA = 1'b0;
            //BOTTOM LEFT 0 COL 0 Row 3
            15'b11010110_0011_000: DATA = 1'b1;
            15'b11010110_0011_001: DATA = 1'b0;
            15'b11010110_0011_010: DATA = 1'b0;
            15'b11010110_0011_011: DATA = 1'b0;
            15'b11010110_0011_100: DATA = 1'b0;
            15'b11010110_0011_101: DATA = 1'b0;
            15'b11010110_0011_110: DATA = 1'b0;
            15'b11010110_0011_111: DATA = 1'b0;
            //BOTTOM LEFT 0 COL 0 Row 4
            15'b11010110_0100_000: DATA = 1'b1;
            15'b11010110_0100_001: DATA = 1'b0;
            15'b11010110_0100_010: DATA = 1'b0;
            15'b11010110_0100_011: DATA = 1'b0;
            15'b11010110_0100_100: DATA = 1'b0;
            15'b11010110_0100_101: DATA = 1'b0;
            15'b11010110_0100_110: DATA = 1'b0;
            15'b11010110_0100_111: DATA = 1'b0;
            //BOTTOM LEFT 0 COL 0 Row 5
            15'b11010110_0101_000: DATA = 1'b1;
            15'b11010110_0101_001: DATA = 1'b0;
            15'b11010110_0101_010: DATA = 1'b0;
            15'b11010110_0101_011: DATA = 1'b0;
            15'b11010110_0101_100: DATA = 1'b0;
            15'b11010110_0101_101: DATA = 1'b0;
            15'b11010110_0101_110: DATA = 1'b0;
            15'b11010110_0101_111: DATA = 1'b0;
            //BOTTOM LEFT 0 COL 0 Row 6
            15'b11010110_0110_000: DATA = 1'b1;
            15'b11010110_0110_001: DATA = 1'b0;
            15'b11010110_0110_010: DATA = 1'b0;
            15'b11010110_0110_011: DATA = 1'b0;
            15'b11010110_0110_100: DATA = 1'b0;
            15'b11010110_0110_101: DATA = 1'b0;
            15'b11010110_0110_110: DATA = 1'b0;
            15'b11010110_0110_111: DATA = 1'b0;
            //BOTTOM LEFT 0 COL 0 Row 7
            15'b11010110_0111_000: DATA = 1'b1;
            15'b11010110_0111_001: DATA = 1'b0;
            15'b11010110_0111_010: DATA = 1'b0;
            15'b11010110_0111_011: DATA = 1'b0;
            15'b11010110_0111_100: DATA = 1'b0;
            15'b11010110_0111_101: DATA = 1'b0;
            15'b11010110_0111_110: DATA = 1'b0;
            15'b11010110_0111_111: DATA = 1'b0;
            //BOTTOM LEFT 0 COL 0 Row 8
            15'b11010110_1000_000: DATA = 1'b1;
            15'b11010110_1000_001: DATA = 1'b0;
            15'b11010110_1000_010: DATA = 1'b0;
            15'b11010110_1000_011: DATA = 1'b0;
            15'b11010110_1000_100: DATA = 1'b0;
            15'b11010110_1000_101: DATA = 1'b0;
            15'b11010110_1000_110: DATA = 1'b0;
            15'b11010110_1000_111: DATA = 1'b0;
            //BOTTOM LEFT 0 COL 0 Row 9
            15'b11010110_1001_000: DATA = 1'b1;
            15'b11010110_1001_001: DATA = 1'b0;
            15'b11010110_1001_010: DATA = 1'b0;
            15'b11010110_1001_011: DATA = 1'b0;
            15'b11010110_1001_100: DATA = 1'b0;
            15'b11010110_1001_101: DATA = 1'b0;
            15'b11010110_1001_110: DATA = 1'b0;
            15'b11010110_1001_111: DATA = 1'b0;
            //BOTTOM LEFT 0 COL 0 Row 10
            15'b11010110_1010_000: DATA = 1'b1;
            15'b11010110_1010_001: DATA = 1'b0;
            15'b11010110_1010_010: DATA = 1'b0;
            15'b11010110_1010_011: DATA = 1'b0;
            15'b11010110_1010_100: DATA = 1'b0;
            15'b11010110_1010_101: DATA = 1'b0;
            15'b11010110_1010_110: DATA = 1'b0;
            15'b11010110_1010_111: DATA = 1'b0;
            //BOTTOM LEFT 0 COL 0 Row 11
            15'b11010110_1011_000: DATA = 1'b1;
            15'b11010110_1011_001: DATA = 1'b0;
            15'b11010110_1011_010: DATA = 1'b0;
            15'b11010110_1011_011: DATA = 1'b0;
            15'b11010110_1011_100: DATA = 1'b0;
            15'b11010110_1011_101: DATA = 1'b0;
            15'b11010110_1011_110: DATA = 1'b0;
            15'b11010110_1011_111: DATA = 1'b0;
            //BOTTOM LEFT 0 COL 0 Row 12
            15'b11010110_1100_000: DATA = 1'b1;
            15'b11010110_1100_001: DATA = 1'b0;
            15'b11010110_1100_010: DATA = 1'b0;
            15'b11010110_1100_011: DATA = 1'b0;
            15'b11010110_1100_100: DATA = 1'b0;
            15'b11010110_1100_101: DATA = 1'b0;
            15'b11010110_1100_110: DATA = 1'b0;
            15'b11010110_1100_111: DATA = 1'b0;
            //BOTTOM LEFT 0 COL 0 Row 13
            15'b11010110_1101_000: DATA = 1'b1;
            15'b11010110_1101_001: DATA = 1'b0;
            15'b11010110_1101_010: DATA = 1'b0;
            15'b11010110_1101_011: DATA = 1'b0;
            15'b11010110_1101_100: DATA = 1'b0;
            15'b11010110_1101_101: DATA = 1'b0;
            15'b11010110_1101_110: DATA = 1'b0;
            15'b11010110_1101_111: DATA = 1'b0;
            //BOTTOM LEFT 0 COL 0 Row 14
            15'b11010110_1110_000: DATA = 1'b1;
            15'b11010110_1110_001: DATA = 1'b0;
            15'b11010110_1110_010: DATA = 1'b0;
            15'b11010110_1110_011: DATA = 1'b0;
            15'b11010110_1110_100: DATA = 1'b0;
            15'b11010110_1110_101: DATA = 1'b0;
            15'b11010110_1110_110: DATA = 1'b0;
            15'b11010110_1110_111: DATA = 1'b0;
            //BOTTOM LEFT 0 COL 0 Row 15
            15'b11010110_1111_000: DATA = 1'b1;
            15'b11010110_1111_001: DATA = 1'b1;
            15'b11010110_1111_010: DATA = 1'b1;
            15'b11010110_1111_011: DATA = 1'b1;
            15'b11010110_1111_100: DATA = 1'b1;
            15'b11010110_1111_101: DATA = 1'b1;
            15'b11010110_1111_110: DATA = 1'b1;
            15'b11010110_1111_111: DATA = 1'b1;
            //BOTTOM RIGHT 0 COL 0 Row 0
            15'b11010111_0000_000: DATA = 1'b0;
            15'b11010111_0000_001: DATA = 1'b0;
            15'b11010111_0000_010: DATA = 1'b0;
            15'b11010111_0000_011: DATA = 1'b0;
            15'b11010111_0000_100: DATA = 1'b0;
            15'b11010111_0000_101: DATA = 1'b0;
            15'b11010111_0000_110: DATA = 1'b0;
            15'b11010111_0000_111: DATA = 1'b1;
            //BOTTOM RIGHT 0 COL 0 Row 1
            15'b11010111_0001_000: DATA = 1'b0;
            15'b11010111_0001_001: DATA = 1'b0;
            15'b11010111_0001_010: DATA = 1'b0;
            15'b11010111_0001_011: DATA = 1'b0;
            15'b11010111_0001_100: DATA = 1'b0;
            15'b11010111_0001_101: DATA = 1'b0;
            15'b11010111_0001_110: DATA = 1'b0;
            15'b11010111_0001_111: DATA = 1'b1;
            //BOTTOM RIGHT 0 COL 0 Row 2
            15'b11010111_0010_000: DATA = 1'b0;
            15'b11010111_0010_001: DATA = 1'b0;
            15'b11010111_0010_010: DATA = 1'b0;
            15'b11010111_0010_011: DATA = 1'b0;
            15'b11010111_0010_100: DATA = 1'b0;
            15'b11010111_0010_101: DATA = 1'b0;
            15'b11010111_0010_110: DATA = 1'b0;
            15'b11010111_0010_111: DATA = 1'b1;
            //BOTTOM RIGHT 0 COL 0 Row 3
            15'b11010111_0011_000: DATA = 1'b0;
            15'b11010111_0011_001: DATA = 1'b0;
            15'b11010111_0011_010: DATA = 1'b0;
            15'b11010111_0011_011: DATA = 1'b0;
            15'b11010111_0011_100: DATA = 1'b0;
            15'b11010111_0011_101: DATA = 1'b0;
            15'b11010111_0011_110: DATA = 1'b0;
            15'b11010111_0011_111: DATA = 1'b1;
            //BOTTOM RIGHT 0 COL 0 Row 4
            15'b11010111_0100_000: DATA = 1'b0;
            15'b11010111_0100_001: DATA = 1'b0;
            15'b11010111_0100_010: DATA = 1'b0;
            15'b11010111_0100_011: DATA = 1'b0;
            15'b11010111_0100_100: DATA = 1'b0;
            15'b11010111_0100_101: DATA = 1'b0;
            15'b11010111_0100_110: DATA = 1'b0;
            15'b11010111_0100_111: DATA = 1'b1;
            //BOTTOM RIGHT 0 COL 0 Row 5
            15'b11010111_0101_000: DATA = 1'b0;
            15'b11010111_0101_001: DATA = 1'b0;
            15'b11010111_0101_010: DATA = 1'b0;
            15'b11010111_0101_011: DATA = 1'b0;
            15'b11010111_0101_100: DATA = 1'b0;
            15'b11010111_0101_101: DATA = 1'b0;
            15'b11010111_0101_110: DATA = 1'b0;
            15'b11010111_0101_111: DATA = 1'b1;
            //BOTTOM RIGHT 0 COL 0 Row 6
            15'b11010111_0110_000: DATA = 1'b0;
            15'b11010111_0110_001: DATA = 1'b0;
            15'b11010111_0110_010: DATA = 1'b0;
            15'b11010111_0110_011: DATA = 1'b0;
            15'b11010111_0110_100: DATA = 1'b0;
            15'b11010111_0110_101: DATA = 1'b0;
            15'b11010111_0110_110: DATA = 1'b0;
            15'b11010111_0110_111: DATA = 1'b1;
            //BOTTOM RIGHT 0 COL 0 Row 7
            15'b11010111_0111_000: DATA = 1'b0;
            15'b11010111_0111_001: DATA = 1'b0;
            15'b11010111_0111_010: DATA = 1'b0;
            15'b11010111_0111_011: DATA = 1'b0;
            15'b11010111_0111_100: DATA = 1'b0;
            15'b11010111_0111_101: DATA = 1'b0;
            15'b11010111_0111_110: DATA = 1'b0;
            15'b11010111_0111_111: DATA = 1'b1;
            //BOTTOM RIGHT 0 COL 0 Row 8
            15'b11010111_1000_000: DATA = 1'b0;
            15'b11010111_1000_001: DATA = 1'b0;
            15'b11010111_1000_010: DATA = 1'b0;
            15'b11010111_1000_011: DATA = 1'b0;
            15'b11010111_1000_100: DATA = 1'b0;
            15'b11010111_1000_101: DATA = 1'b0;
            15'b11010111_1000_110: DATA = 1'b0;
            15'b11010111_1000_111: DATA = 1'b1;
            //BOTTOM RIGHT 0 COL 0 Row 9
            15'b11010111_1001_000: DATA = 1'b0;
            15'b11010111_1001_001: DATA = 1'b0;
            15'b11010111_1001_010: DATA = 1'b0;
            15'b11010111_1001_011: DATA = 1'b0;
            15'b11010111_1001_100: DATA = 1'b0;
            15'b11010111_1001_101: DATA = 1'b0;
            15'b11010111_1001_110: DATA = 1'b0;
            15'b11010111_1001_111: DATA = 1'b1;
            //BOTTOM RIGHT 0 COL 0 Row 10
            15'b11010111_1010_000: DATA = 1'b0;
            15'b11010111_1010_001: DATA = 1'b0;
            15'b11010111_1010_010: DATA = 1'b0;
            15'b11010111_1010_011: DATA = 1'b0;
            15'b11010111_1010_100: DATA = 1'b0;
            15'b11010111_1010_101: DATA = 1'b0;
            15'b11010111_1010_110: DATA = 1'b0;
            15'b11010111_1010_111: DATA = 1'b1;
            //BOTTOM RIGHT 0 COL 0 Row 11
            15'b11010111_1011_000: DATA = 1'b0;
            15'b11010111_1011_001: DATA = 1'b0;
            15'b11010111_1011_010: DATA = 1'b0;
            15'b11010111_1011_011: DATA = 1'b0;
            15'b11010111_1011_100: DATA = 1'b0;
            15'b11010111_1011_101: DATA = 1'b0;
            15'b11010111_1011_110: DATA = 1'b0;
            15'b11010111_1011_111: DATA = 1'b1;
            //BOTTOM RIGHT 0 COL 0 Row 12
            15'b11010111_1100_000: DATA = 1'b0;
            15'b11010111_1100_001: DATA = 1'b0;
            15'b11010111_1100_010: DATA = 1'b0;
            15'b11010111_1100_011: DATA = 1'b0;
            15'b11010111_1100_100: DATA = 1'b0;
            15'b11010111_1100_101: DATA = 1'b0;
            15'b11010111_1100_110: DATA = 1'b0;
            15'b11010111_1100_111: DATA = 1'b1;
            //BOTTOM RIGHT 0 COL 0 Row 13
            15'b11010111_1101_000: DATA = 1'b0;
            15'b11010111_1101_001: DATA = 1'b0;
            15'b11010111_1101_010: DATA = 1'b0;
            15'b11010111_1101_011: DATA = 1'b0;
            15'b11010111_1101_100: DATA = 1'b0;
            15'b11010111_1101_101: DATA = 1'b0;
            15'b11010111_1101_110: DATA = 1'b0;
            15'b11010111_1101_111: DATA = 1'b1;
            //BOTTOM RIGHT 0 COL 0 Row 14
            15'b11010111_1110_000: DATA = 1'b0;
            15'b11010111_1110_001: DATA = 1'b0;
            15'b11010111_1110_010: DATA = 1'b0;
            15'b11010111_1110_011: DATA = 1'b0;
            15'b11010111_1110_100: DATA = 1'b0;
            15'b11010111_1110_101: DATA = 1'b0;
            15'b11010111_1110_110: DATA = 1'b0;
            15'b11010111_1110_111: DATA = 1'b1;
            //BOTTOM RIGHT 0 COL 0 Row 15
            15'b11010111_1111_000: DATA = 1'b1;
            15'b11010111_1111_001: DATA = 1'b1;
            15'b11010111_1111_010: DATA = 1'b1;
            15'b11010111_1111_011: DATA = 1'b1;
            15'b11010111_1111_100: DATA = 1'b1;
            15'b11010111_1111_101: DATA = 1'b1;
            15'b11010111_1111_110: DATA = 1'b1;
            15'b11010111_1111_111: DATA = 1'b1;
            //SAWTOOTHY+ ROW 0 COL 0 Row 0
            15'b11011000_0000_000: DATA = 1'b1;
            15'b11011000_0000_001: DATA = 1'b1;
            15'b11011000_0000_010: DATA = 1'b0;
            15'b11011000_0000_011: DATA = 1'b0;
            15'b11011000_0000_100: DATA = 1'b0;
            15'b11011000_0000_101: DATA = 1'b0;
            15'b11011000_0000_110: DATA = 1'b0;
            15'b11011000_0000_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 0 Row 1
            15'b11011000_0001_000: DATA = 1'b1;
            15'b11011000_0001_001: DATA = 1'b0;
            15'b11011000_0001_010: DATA = 1'b1;
            15'b11011000_0001_011: DATA = 1'b0;
            15'b11011000_0001_100: DATA = 1'b0;
            15'b11011000_0001_101: DATA = 1'b0;
            15'b11011000_0001_110: DATA = 1'b0;
            15'b11011000_0001_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 0 Row 2
            15'b11011000_0010_000: DATA = 1'b1;
            15'b11011000_0010_001: DATA = 1'b0;
            15'b11011000_0010_010: DATA = 1'b1;
            15'b11011000_0010_011: DATA = 1'b1;
            15'b11011000_0010_100: DATA = 1'b0;
            15'b11011000_0010_101: DATA = 1'b0;
            15'b11011000_0010_110: DATA = 1'b0;
            15'b11011000_0010_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 0 Row 3
            15'b11011000_0011_000: DATA = 1'b1;
            15'b11011000_0011_001: DATA = 1'b0;
            15'b11011000_0011_010: DATA = 1'b0;
            15'b11011000_0011_011: DATA = 1'b1;
            15'b11011000_0011_100: DATA = 1'b1;
            15'b11011000_0011_101: DATA = 1'b0;
            15'b11011000_0011_110: DATA = 1'b0;
            15'b11011000_0011_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 0 Row 4
            15'b11011000_0100_000: DATA = 1'b1;
            15'b11011000_0100_001: DATA = 1'b0;
            15'b11011000_0100_010: DATA = 1'b0;
            15'b11011000_0100_011: DATA = 1'b0;
            15'b11011000_0100_100: DATA = 1'b1;
            15'b11011000_0100_101: DATA = 1'b1;
            15'b11011000_0100_110: DATA = 1'b1;
            15'b11011000_0100_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 0 Row 5
            15'b11011000_0101_000: DATA = 1'b1;
            15'b11011000_0101_001: DATA = 1'b0;
            15'b11011000_0101_010: DATA = 1'b0;
            15'b11011000_0101_011: DATA = 1'b0;
            15'b11011000_0101_100: DATA = 1'b0;
            15'b11011000_0101_101: DATA = 1'b0;
            15'b11011000_0101_110: DATA = 1'b1;
            15'b11011000_0101_111: DATA = 1'b1;
            //SAWTOOTHY+ ROW 0 COL 0 Row 6
            15'b11011000_0110_000: DATA = 1'b1;
            15'b11011000_0110_001: DATA = 1'b0;
            15'b11011000_0110_010: DATA = 1'b0;
            15'b11011000_0110_011: DATA = 1'b0;
            15'b11011000_0110_100: DATA = 1'b0;
            15'b11011000_0110_101: DATA = 1'b0;
            15'b11011000_0110_110: DATA = 1'b0;
            15'b11011000_0110_111: DATA = 1'b1;
            //SAWTOOTHY+ ROW 0 COL 0 Row 7
            15'b11011000_0111_000: DATA = 1'b1;
            15'b11011000_0111_001: DATA = 1'b0;
            15'b11011000_0111_010: DATA = 1'b0;
            15'b11011000_0111_011: DATA = 1'b0;
            15'b11011000_0111_100: DATA = 1'b0;
            15'b11011000_0111_101: DATA = 1'b0;
            15'b11011000_0111_110: DATA = 1'b0;
            15'b11011000_0111_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 0 Row 8
            15'b11011000_1000_000: DATA = 1'b1;
            15'b11011000_1000_001: DATA = 1'b0;
            15'b11011000_1000_010: DATA = 1'b0;
            15'b11011000_1000_011: DATA = 1'b0;
            15'b11011000_1000_100: DATA = 1'b0;
            15'b11011000_1000_101: DATA = 1'b0;
            15'b11011000_1000_110: DATA = 1'b0;
            15'b11011000_1000_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 0 Row 9
            15'b11011000_1001_000: DATA = 1'b1;
            15'b11011000_1001_001: DATA = 1'b0;
            15'b11011000_1001_010: DATA = 1'b0;
            15'b11011000_1001_011: DATA = 1'b0;
            15'b11011000_1001_100: DATA = 1'b0;
            15'b11011000_1001_101: DATA = 1'b0;
            15'b11011000_1001_110: DATA = 1'b0;
            15'b11011000_1001_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 0 Row 10
            15'b11011000_1010_000: DATA = 1'b1;
            15'b11011000_1010_001: DATA = 1'b0;
            15'b11011000_1010_010: DATA = 1'b0;
            15'b11011000_1010_011: DATA = 1'b0;
            15'b11011000_1010_100: DATA = 1'b0;
            15'b11011000_1010_101: DATA = 1'b0;
            15'b11011000_1010_110: DATA = 1'b0;
            15'b11011000_1010_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 0 Row 11
            15'b11011000_1011_000: DATA = 1'b1;
            15'b11011000_1011_001: DATA = 1'b0;
            15'b11011000_1011_010: DATA = 1'b0;
            15'b11011000_1011_011: DATA = 1'b0;
            15'b11011000_1011_100: DATA = 1'b0;
            15'b11011000_1011_101: DATA = 1'b0;
            15'b11011000_1011_110: DATA = 1'b0;
            15'b11011000_1011_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 0 Row 12
            15'b11011000_1100_000: DATA = 1'b1;
            15'b11011000_1100_001: DATA = 1'b0;
            15'b11011000_1100_010: DATA = 1'b0;
            15'b11011000_1100_011: DATA = 1'b0;
            15'b11011000_1100_100: DATA = 1'b0;
            15'b11011000_1100_101: DATA = 1'b0;
            15'b11011000_1100_110: DATA = 1'b0;
            15'b11011000_1100_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 0 Row 13
            15'b11011000_1101_000: DATA = 1'b1;
            15'b11011000_1101_001: DATA = 1'b0;
            15'b11011000_1101_010: DATA = 1'b0;
            15'b11011000_1101_011: DATA = 1'b0;
            15'b11011000_1101_100: DATA = 1'b0;
            15'b11011000_1101_101: DATA = 1'b0;
            15'b11011000_1101_110: DATA = 1'b0;
            15'b11011000_1101_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 0 Row 14
            15'b11011000_1110_000: DATA = 1'b1;
            15'b11011000_1110_001: DATA = 1'b0;
            15'b11011000_1110_010: DATA = 1'b0;
            15'b11011000_1110_011: DATA = 1'b0;
            15'b11011000_1110_100: DATA = 1'b0;
            15'b11011000_1110_101: DATA = 1'b0;
            15'b11011000_1110_110: DATA = 1'b0;
            15'b11011000_1110_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 0 Row 15
            15'b11011000_1111_000: DATA = 1'b1;
            15'b11011000_1111_001: DATA = 1'b0;
            15'b11011000_1111_010: DATA = 1'b0;
            15'b11011000_1111_011: DATA = 1'b0;
            15'b11011000_1111_100: DATA = 1'b0;
            15'b11011000_1111_101: DATA = 1'b0;
            15'b11011000_1111_110: DATA = 1'b0;
            15'b11011000_1111_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 1 Row 0
            15'b11011001_0000_000: DATA = 1'b0;
            15'b11011001_0000_001: DATA = 1'b0;
            15'b11011001_0000_010: DATA = 1'b0;
            15'b11011001_0000_011: DATA = 1'b0;
            15'b11011001_0000_100: DATA = 1'b0;
            15'b11011001_0000_101: DATA = 1'b0;
            15'b11011001_0000_110: DATA = 1'b0;
            15'b11011001_0000_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 1 Row 1
            15'b11011001_0001_000: DATA = 1'b0;
            15'b11011001_0001_001: DATA = 1'b0;
            15'b11011001_0001_010: DATA = 1'b0;
            15'b11011001_0001_011: DATA = 1'b0;
            15'b11011001_0001_100: DATA = 1'b0;
            15'b11011001_0001_101: DATA = 1'b0;
            15'b11011001_0001_110: DATA = 1'b0;
            15'b11011001_0001_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 1 Row 2
            15'b11011001_0010_000: DATA = 1'b0;
            15'b11011001_0010_001: DATA = 1'b0;
            15'b11011001_0010_010: DATA = 1'b0;
            15'b11011001_0010_011: DATA = 1'b0;
            15'b11011001_0010_100: DATA = 1'b0;
            15'b11011001_0010_101: DATA = 1'b0;
            15'b11011001_0010_110: DATA = 1'b0;
            15'b11011001_0010_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 1 Row 3
            15'b11011001_0011_000: DATA = 1'b0;
            15'b11011001_0011_001: DATA = 1'b0;
            15'b11011001_0011_010: DATA = 1'b0;
            15'b11011001_0011_011: DATA = 1'b0;
            15'b11011001_0011_100: DATA = 1'b0;
            15'b11011001_0011_101: DATA = 1'b0;
            15'b11011001_0011_110: DATA = 1'b0;
            15'b11011001_0011_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 1 Row 4
            15'b11011001_0100_000: DATA = 1'b0;
            15'b11011001_0100_001: DATA = 1'b0;
            15'b11011001_0100_010: DATA = 1'b0;
            15'b11011001_0100_011: DATA = 1'b0;
            15'b11011001_0100_100: DATA = 1'b0;
            15'b11011001_0100_101: DATA = 1'b0;
            15'b11011001_0100_110: DATA = 1'b0;
            15'b11011001_0100_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 1 Row 5
            15'b11011001_0101_000: DATA = 1'b0;
            15'b11011001_0101_001: DATA = 1'b0;
            15'b11011001_0101_010: DATA = 1'b0;
            15'b11011001_0101_011: DATA = 1'b0;
            15'b11011001_0101_100: DATA = 1'b0;
            15'b11011001_0101_101: DATA = 1'b0;
            15'b11011001_0101_110: DATA = 1'b0;
            15'b11011001_0101_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 1 Row 6
            15'b11011001_0110_000: DATA = 1'b1;
            15'b11011001_0110_001: DATA = 1'b0;
            15'b11011001_0110_010: DATA = 1'b0;
            15'b11011001_0110_011: DATA = 1'b0;
            15'b11011001_0110_100: DATA = 1'b0;
            15'b11011001_0110_101: DATA = 1'b0;
            15'b11011001_0110_110: DATA = 1'b0;
            15'b11011001_0110_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 1 Row 7
            15'b11011001_0111_000: DATA = 1'b1;
            15'b11011001_0111_001: DATA = 1'b1;
            15'b11011001_0111_010: DATA = 1'b0;
            15'b11011001_0111_011: DATA = 1'b0;
            15'b11011001_0111_100: DATA = 1'b0;
            15'b11011001_0111_101: DATA = 1'b0;
            15'b11011001_0111_110: DATA = 1'b0;
            15'b11011001_0111_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 1 Row 8
            15'b11011001_1000_000: DATA = 1'b0;
            15'b11011001_1000_001: DATA = 1'b1;
            15'b11011001_1000_010: DATA = 1'b1;
            15'b11011001_1000_011: DATA = 1'b1;
            15'b11011001_1000_100: DATA = 1'b0;
            15'b11011001_1000_101: DATA = 1'b0;
            15'b11011001_1000_110: DATA = 1'b0;
            15'b11011001_1000_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 1 Row 9
            15'b11011001_1001_000: DATA = 1'b0;
            15'b11011001_1001_001: DATA = 1'b0;
            15'b11011001_1001_010: DATA = 1'b0;
            15'b11011001_1001_011: DATA = 1'b1;
            15'b11011001_1001_100: DATA = 1'b1;
            15'b11011001_1001_101: DATA = 1'b0;
            15'b11011001_1001_110: DATA = 1'b0;
            15'b11011001_1001_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 1 Row 10
            15'b11011001_1010_000: DATA = 1'b0;
            15'b11011001_1010_001: DATA = 1'b0;
            15'b11011001_1010_010: DATA = 1'b0;
            15'b11011001_1010_011: DATA = 1'b0;
            15'b11011001_1010_100: DATA = 1'b1;
            15'b11011001_1010_101: DATA = 1'b1;
            15'b11011001_1010_110: DATA = 1'b0;
            15'b11011001_1010_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 1 Row 11
            15'b11011001_1011_000: DATA = 1'b0;
            15'b11011001_1011_001: DATA = 1'b0;
            15'b11011001_1011_010: DATA = 1'b0;
            15'b11011001_1011_011: DATA = 1'b0;
            15'b11011001_1011_100: DATA = 1'b0;
            15'b11011001_1011_101: DATA = 1'b1;
            15'b11011001_1011_110: DATA = 1'b1;
            15'b11011001_1011_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 1 Row 12
            15'b11011001_1100_000: DATA = 1'b0;
            15'b11011001_1100_001: DATA = 1'b0;
            15'b11011001_1100_010: DATA = 1'b0;
            15'b11011001_1100_011: DATA = 1'b0;
            15'b11011001_1100_100: DATA = 1'b0;
            15'b11011001_1100_101: DATA = 1'b0;
            15'b11011001_1100_110: DATA = 1'b1;
            15'b11011001_1100_111: DATA = 1'b1;
            //SAWTOOTHY+ ROW 0 COL 1 Row 13
            15'b11011001_1101_000: DATA = 1'b0;
            15'b11011001_1101_001: DATA = 1'b0;
            15'b11011001_1101_010: DATA = 1'b0;
            15'b11011001_1101_011: DATA = 1'b0;
            15'b11011001_1101_100: DATA = 1'b0;
            15'b11011001_1101_101: DATA = 1'b0;
            15'b11011001_1101_110: DATA = 1'b0;
            15'b11011001_1101_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 1 Row 14
            15'b11011001_1110_000: DATA = 1'b0;
            15'b11011001_1110_001: DATA = 1'b0;
            15'b11011001_1110_010: DATA = 1'b0;
            15'b11011001_1110_011: DATA = 1'b0;
            15'b11011001_1110_100: DATA = 1'b0;
            15'b11011001_1110_101: DATA = 1'b0;
            15'b11011001_1110_110: DATA = 1'b0;
            15'b11011001_1110_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 1 Row 15
            15'b11011001_1111_000: DATA = 1'b0;
            15'b11011001_1111_001: DATA = 1'b0;
            15'b11011001_1111_010: DATA = 1'b0;
            15'b11011001_1111_011: DATA = 1'b0;
            15'b11011001_1111_100: DATA = 1'b0;
            15'b11011001_1111_101: DATA = 1'b0;
            15'b11011001_1111_110: DATA = 1'b0;
            15'b11011001_1111_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 2 Row 0
            15'b11011010_0000_000: DATA = 1'b0;
            15'b11011010_0000_001: DATA = 1'b0;
            15'b11011010_0000_010: DATA = 1'b0;
            15'b11011010_0000_011: DATA = 1'b0;
            15'b11011010_0000_100: DATA = 1'b0;
            15'b11011010_0000_101: DATA = 1'b0;
            15'b11011010_0000_110: DATA = 1'b0;
            15'b11011010_0000_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 2 Row 1
            15'b11011010_0001_000: DATA = 1'b0;
            15'b11011010_0001_001: DATA = 1'b0;
            15'b11011010_0001_010: DATA = 1'b0;
            15'b11011010_0001_011: DATA = 1'b0;
            15'b11011010_0001_100: DATA = 1'b0;
            15'b11011010_0001_101: DATA = 1'b0;
            15'b11011010_0001_110: DATA = 1'b0;
            15'b11011010_0001_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 2 Row 2
            15'b11011010_0010_000: DATA = 1'b0;
            15'b11011010_0010_001: DATA = 1'b0;
            15'b11011010_0010_010: DATA = 1'b0;
            15'b11011010_0010_011: DATA = 1'b0;
            15'b11011010_0010_100: DATA = 1'b0;
            15'b11011010_0010_101: DATA = 1'b0;
            15'b11011010_0010_110: DATA = 1'b0;
            15'b11011010_0010_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 2 Row 3
            15'b11011010_0011_000: DATA = 1'b0;
            15'b11011010_0011_001: DATA = 1'b0;
            15'b11011010_0011_010: DATA = 1'b0;
            15'b11011010_0011_011: DATA = 1'b0;
            15'b11011010_0011_100: DATA = 1'b0;
            15'b11011010_0011_101: DATA = 1'b0;
            15'b11011010_0011_110: DATA = 1'b0;
            15'b11011010_0011_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 2 Row 4
            15'b11011010_0100_000: DATA = 1'b0;
            15'b11011010_0100_001: DATA = 1'b0;
            15'b11011010_0100_010: DATA = 1'b0;
            15'b11011010_0100_011: DATA = 1'b0;
            15'b11011010_0100_100: DATA = 1'b0;
            15'b11011010_0100_101: DATA = 1'b0;
            15'b11011010_0100_110: DATA = 1'b0;
            15'b11011010_0100_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 2 Row 5
            15'b11011010_0101_000: DATA = 1'b0;
            15'b11011010_0101_001: DATA = 1'b0;
            15'b11011010_0101_010: DATA = 1'b0;
            15'b11011010_0101_011: DATA = 1'b0;
            15'b11011010_0101_100: DATA = 1'b0;
            15'b11011010_0101_101: DATA = 1'b0;
            15'b11011010_0101_110: DATA = 1'b0;
            15'b11011010_0101_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 2 Row 6
            15'b11011010_0110_000: DATA = 1'b0;
            15'b11011010_0110_001: DATA = 1'b0;
            15'b11011010_0110_010: DATA = 1'b0;
            15'b11011010_0110_011: DATA = 1'b0;
            15'b11011010_0110_100: DATA = 1'b0;
            15'b11011010_0110_101: DATA = 1'b0;
            15'b11011010_0110_110: DATA = 1'b0;
            15'b11011010_0110_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 2 Row 7
            15'b11011010_0111_000: DATA = 1'b0;
            15'b11011010_0111_001: DATA = 1'b0;
            15'b11011010_0111_010: DATA = 1'b0;
            15'b11011010_0111_011: DATA = 1'b0;
            15'b11011010_0111_100: DATA = 1'b0;
            15'b11011010_0111_101: DATA = 1'b0;
            15'b11011010_0111_110: DATA = 1'b0;
            15'b11011010_0111_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 2 Row 8
            15'b11011010_1000_000: DATA = 1'b0;
            15'b11011010_1000_001: DATA = 1'b0;
            15'b11011010_1000_010: DATA = 1'b0;
            15'b11011010_1000_011: DATA = 1'b0;
            15'b11011010_1000_100: DATA = 1'b0;
            15'b11011010_1000_101: DATA = 1'b0;
            15'b11011010_1000_110: DATA = 1'b0;
            15'b11011010_1000_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 2 Row 9
            15'b11011010_1001_000: DATA = 1'b0;
            15'b11011010_1001_001: DATA = 1'b0;
            15'b11011010_1001_010: DATA = 1'b0;
            15'b11011010_1001_011: DATA = 1'b0;
            15'b11011010_1001_100: DATA = 1'b0;
            15'b11011010_1001_101: DATA = 1'b0;
            15'b11011010_1001_110: DATA = 1'b0;
            15'b11011010_1001_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 2 Row 10
            15'b11011010_1010_000: DATA = 1'b0;
            15'b11011010_1010_001: DATA = 1'b0;
            15'b11011010_1010_010: DATA = 1'b0;
            15'b11011010_1010_011: DATA = 1'b0;
            15'b11011010_1010_100: DATA = 1'b0;
            15'b11011010_1010_101: DATA = 1'b0;
            15'b11011010_1010_110: DATA = 1'b0;
            15'b11011010_1010_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 2 Row 11
            15'b11011010_1011_000: DATA = 1'b0;
            15'b11011010_1011_001: DATA = 1'b0;
            15'b11011010_1011_010: DATA = 1'b0;
            15'b11011010_1011_011: DATA = 1'b0;
            15'b11011010_1011_100: DATA = 1'b0;
            15'b11011010_1011_101: DATA = 1'b0;
            15'b11011010_1011_110: DATA = 1'b0;
            15'b11011010_1011_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 2 Row 12
            15'b11011010_1100_000: DATA = 1'b1;
            15'b11011010_1100_001: DATA = 1'b0;
            15'b11011010_1100_010: DATA = 1'b0;
            15'b11011010_1100_011: DATA = 1'b0;
            15'b11011010_1100_100: DATA = 1'b0;
            15'b11011010_1100_101: DATA = 1'b0;
            15'b11011010_1100_110: DATA = 1'b0;
            15'b11011010_1100_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 2 Row 13
            15'b11011010_1101_000: DATA = 1'b1;
            15'b11011010_1101_001: DATA = 1'b1;
            15'b11011010_1101_010: DATA = 1'b0;
            15'b11011010_1101_011: DATA = 1'b0;
            15'b11011010_1101_100: DATA = 1'b0;
            15'b11011010_1101_101: DATA = 1'b0;
            15'b11011010_1101_110: DATA = 1'b0;
            15'b11011010_1101_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 2 Row 14
            15'b11011010_1110_000: DATA = 1'b0;
            15'b11011010_1110_001: DATA = 1'b1;
            15'b11011010_1110_010: DATA = 1'b1;
            15'b11011010_1110_011: DATA = 1'b0;
            15'b11011010_1110_100: DATA = 1'b0;
            15'b11011010_1110_101: DATA = 1'b0;
            15'b11011010_1110_110: DATA = 1'b0;
            15'b11011010_1110_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 2 Row 15
            15'b11011010_1111_000: DATA = 1'b0;
            15'b11011010_1111_001: DATA = 1'b0;
            15'b11011010_1111_010: DATA = 1'b1;
            15'b11011010_1111_011: DATA = 1'b1;
            15'b11011010_1111_100: DATA = 1'b0;
            15'b11011010_1111_101: DATA = 1'b0;
            15'b11011010_1111_110: DATA = 1'b0;
            15'b11011010_1111_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 3 Row 0
            15'b11011011_0000_000: DATA = 1'b0;
            15'b11011011_0000_001: DATA = 1'b0;
            15'b11011011_0000_010: DATA = 1'b0;
            15'b11011011_0000_011: DATA = 1'b0;
            15'b11011011_0000_100: DATA = 1'b0;
            15'b11011011_0000_101: DATA = 1'b0;
            15'b11011011_0000_110: DATA = 1'b0;
            15'b11011011_0000_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 3 Row 1
            15'b11011011_0001_000: DATA = 1'b0;
            15'b11011011_0001_001: DATA = 1'b0;
            15'b11011011_0001_010: DATA = 1'b0;
            15'b11011011_0001_011: DATA = 1'b0;
            15'b11011011_0001_100: DATA = 1'b0;
            15'b11011011_0001_101: DATA = 1'b0;
            15'b11011011_0001_110: DATA = 1'b0;
            15'b11011011_0001_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 3 Row 2
            15'b11011011_0010_000: DATA = 1'b0;
            15'b11011011_0010_001: DATA = 1'b0;
            15'b11011011_0010_010: DATA = 1'b0;
            15'b11011011_0010_011: DATA = 1'b0;
            15'b11011011_0010_100: DATA = 1'b0;
            15'b11011011_0010_101: DATA = 1'b0;
            15'b11011011_0010_110: DATA = 1'b0;
            15'b11011011_0010_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 3 Row 3
            15'b11011011_0011_000: DATA = 1'b0;
            15'b11011011_0011_001: DATA = 1'b0;
            15'b11011011_0011_010: DATA = 1'b0;
            15'b11011011_0011_011: DATA = 1'b0;
            15'b11011011_0011_100: DATA = 1'b0;
            15'b11011011_0011_101: DATA = 1'b0;
            15'b11011011_0011_110: DATA = 1'b0;
            15'b11011011_0011_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 3 Row 4
            15'b11011011_0100_000: DATA = 1'b0;
            15'b11011011_0100_001: DATA = 1'b0;
            15'b11011011_0100_010: DATA = 1'b0;
            15'b11011011_0100_011: DATA = 1'b0;
            15'b11011011_0100_100: DATA = 1'b0;
            15'b11011011_0100_101: DATA = 1'b0;
            15'b11011011_0100_110: DATA = 1'b0;
            15'b11011011_0100_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 3 Row 5
            15'b11011011_0101_000: DATA = 1'b0;
            15'b11011011_0101_001: DATA = 1'b0;
            15'b11011011_0101_010: DATA = 1'b0;
            15'b11011011_0101_011: DATA = 1'b0;
            15'b11011011_0101_100: DATA = 1'b0;
            15'b11011011_0101_101: DATA = 1'b0;
            15'b11011011_0101_110: DATA = 1'b0;
            15'b11011011_0101_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 3 Row 6
            15'b11011011_0110_000: DATA = 1'b0;
            15'b11011011_0110_001: DATA = 1'b0;
            15'b11011011_0110_010: DATA = 1'b0;
            15'b11011011_0110_011: DATA = 1'b0;
            15'b11011011_0110_100: DATA = 1'b0;
            15'b11011011_0110_101: DATA = 1'b0;
            15'b11011011_0110_110: DATA = 1'b0;
            15'b11011011_0110_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 3 Row 7
            15'b11011011_0111_000: DATA = 1'b0;
            15'b11011011_0111_001: DATA = 1'b0;
            15'b11011011_0111_010: DATA = 1'b0;
            15'b11011011_0111_011: DATA = 1'b0;
            15'b11011011_0111_100: DATA = 1'b0;
            15'b11011011_0111_101: DATA = 1'b0;
            15'b11011011_0111_110: DATA = 1'b0;
            15'b11011011_0111_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 3 Row 8
            15'b11011011_1000_000: DATA = 1'b0;
            15'b11011011_1000_001: DATA = 1'b0;
            15'b11011011_1000_010: DATA = 1'b0;
            15'b11011011_1000_011: DATA = 1'b0;
            15'b11011011_1000_100: DATA = 1'b0;
            15'b11011011_1000_101: DATA = 1'b0;
            15'b11011011_1000_110: DATA = 1'b0;
            15'b11011011_1000_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 3 Row 9
            15'b11011011_1001_000: DATA = 1'b0;
            15'b11011011_1001_001: DATA = 1'b0;
            15'b11011011_1001_010: DATA = 1'b0;
            15'b11011011_1001_011: DATA = 1'b0;
            15'b11011011_1001_100: DATA = 1'b0;
            15'b11011011_1001_101: DATA = 1'b0;
            15'b11011011_1001_110: DATA = 1'b0;
            15'b11011011_1001_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 3 Row 10
            15'b11011011_1010_000: DATA = 1'b0;
            15'b11011011_1010_001: DATA = 1'b0;
            15'b11011011_1010_010: DATA = 1'b0;
            15'b11011011_1010_011: DATA = 1'b0;
            15'b11011011_1010_100: DATA = 1'b0;
            15'b11011011_1010_101: DATA = 1'b0;
            15'b11011011_1010_110: DATA = 1'b0;
            15'b11011011_1010_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 3 Row 11
            15'b11011011_1011_000: DATA = 1'b0;
            15'b11011011_1011_001: DATA = 1'b0;
            15'b11011011_1011_010: DATA = 1'b0;
            15'b11011011_1011_011: DATA = 1'b0;
            15'b11011011_1011_100: DATA = 1'b0;
            15'b11011011_1011_101: DATA = 1'b0;
            15'b11011011_1011_110: DATA = 1'b0;
            15'b11011011_1011_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 3 Row 12
            15'b11011011_1100_000: DATA = 1'b0;
            15'b11011011_1100_001: DATA = 1'b0;
            15'b11011011_1100_010: DATA = 1'b0;
            15'b11011011_1100_011: DATA = 1'b0;
            15'b11011011_1100_100: DATA = 1'b0;
            15'b11011011_1100_101: DATA = 1'b0;
            15'b11011011_1100_110: DATA = 1'b0;
            15'b11011011_1100_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 3 Row 13
            15'b11011011_1101_000: DATA = 1'b0;
            15'b11011011_1101_001: DATA = 1'b0;
            15'b11011011_1101_010: DATA = 1'b0;
            15'b11011011_1101_011: DATA = 1'b0;
            15'b11011011_1101_100: DATA = 1'b0;
            15'b11011011_1101_101: DATA = 1'b0;
            15'b11011011_1101_110: DATA = 1'b0;
            15'b11011011_1101_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 3 Row 14
            15'b11011011_1110_000: DATA = 1'b0;
            15'b11011011_1110_001: DATA = 1'b0;
            15'b11011011_1110_010: DATA = 1'b0;
            15'b11011011_1110_011: DATA = 1'b0;
            15'b11011011_1110_100: DATA = 1'b0;
            15'b11011011_1110_101: DATA = 1'b0;
            15'b11011011_1110_110: DATA = 1'b0;
            15'b11011011_1110_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 3 Row 15
            15'b11011011_1111_000: DATA = 1'b0;
            15'b11011011_1111_001: DATA = 1'b0;
            15'b11011011_1111_010: DATA = 1'b0;
            15'b11011011_1111_011: DATA = 1'b0;
            15'b11011011_1111_100: DATA = 1'b0;
            15'b11011011_1111_101: DATA = 1'b0;
            15'b11011011_1111_110: DATA = 1'b0;
            15'b11011011_1111_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 4 Row 0
            15'b11011100_0000_000: DATA = 1'b0;
            15'b11011100_0000_001: DATA = 1'b0;
            15'b11011100_0000_010: DATA = 1'b0;
            15'b11011100_0000_011: DATA = 1'b0;
            15'b11011100_0000_100: DATA = 1'b0;
            15'b11011100_0000_101: DATA = 1'b0;
            15'b11011100_0000_110: DATA = 1'b0;
            15'b11011100_0000_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 4 Row 1
            15'b11011100_0001_000: DATA = 1'b0;
            15'b11011100_0001_001: DATA = 1'b0;
            15'b11011100_0001_010: DATA = 1'b0;
            15'b11011100_0001_011: DATA = 1'b0;
            15'b11011100_0001_100: DATA = 1'b0;
            15'b11011100_0001_101: DATA = 1'b0;
            15'b11011100_0001_110: DATA = 1'b0;
            15'b11011100_0001_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 4 Row 2
            15'b11011100_0010_000: DATA = 1'b0;
            15'b11011100_0010_001: DATA = 1'b0;
            15'b11011100_0010_010: DATA = 1'b0;
            15'b11011100_0010_011: DATA = 1'b0;
            15'b11011100_0010_100: DATA = 1'b0;
            15'b11011100_0010_101: DATA = 1'b0;
            15'b11011100_0010_110: DATA = 1'b0;
            15'b11011100_0010_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 4 Row 3
            15'b11011100_0011_000: DATA = 1'b0;
            15'b11011100_0011_001: DATA = 1'b0;
            15'b11011100_0011_010: DATA = 1'b0;
            15'b11011100_0011_011: DATA = 1'b0;
            15'b11011100_0011_100: DATA = 1'b0;
            15'b11011100_0011_101: DATA = 1'b0;
            15'b11011100_0011_110: DATA = 1'b0;
            15'b11011100_0011_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 4 Row 4
            15'b11011100_0100_000: DATA = 1'b0;
            15'b11011100_0100_001: DATA = 1'b0;
            15'b11011100_0100_010: DATA = 1'b0;
            15'b11011100_0100_011: DATA = 1'b0;
            15'b11011100_0100_100: DATA = 1'b0;
            15'b11011100_0100_101: DATA = 1'b0;
            15'b11011100_0100_110: DATA = 1'b0;
            15'b11011100_0100_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 4 Row 5
            15'b11011100_0101_000: DATA = 1'b0;
            15'b11011100_0101_001: DATA = 1'b0;
            15'b11011100_0101_010: DATA = 1'b0;
            15'b11011100_0101_011: DATA = 1'b0;
            15'b11011100_0101_100: DATA = 1'b0;
            15'b11011100_0101_101: DATA = 1'b0;
            15'b11011100_0101_110: DATA = 1'b0;
            15'b11011100_0101_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 4 Row 6
            15'b11011100_0110_000: DATA = 1'b0;
            15'b11011100_0110_001: DATA = 1'b0;
            15'b11011100_0110_010: DATA = 1'b0;
            15'b11011100_0110_011: DATA = 1'b0;
            15'b11011100_0110_100: DATA = 1'b0;
            15'b11011100_0110_101: DATA = 1'b0;
            15'b11011100_0110_110: DATA = 1'b0;
            15'b11011100_0110_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 4 Row 7
            15'b11011100_0111_000: DATA = 1'b0;
            15'b11011100_0111_001: DATA = 1'b0;
            15'b11011100_0111_010: DATA = 1'b0;
            15'b11011100_0111_011: DATA = 1'b0;
            15'b11011100_0111_100: DATA = 1'b0;
            15'b11011100_0111_101: DATA = 1'b0;
            15'b11011100_0111_110: DATA = 1'b0;
            15'b11011100_0111_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 4 Row 8
            15'b11011100_1000_000: DATA = 1'b0;
            15'b11011100_1000_001: DATA = 1'b0;
            15'b11011100_1000_010: DATA = 1'b0;
            15'b11011100_1000_011: DATA = 1'b0;
            15'b11011100_1000_100: DATA = 1'b0;
            15'b11011100_1000_101: DATA = 1'b0;
            15'b11011100_1000_110: DATA = 1'b0;
            15'b11011100_1000_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 4 Row 9
            15'b11011100_1001_000: DATA = 1'b0;
            15'b11011100_1001_001: DATA = 1'b0;
            15'b11011100_1001_010: DATA = 1'b0;
            15'b11011100_1001_011: DATA = 1'b0;
            15'b11011100_1001_100: DATA = 1'b0;
            15'b11011100_1001_101: DATA = 1'b0;
            15'b11011100_1001_110: DATA = 1'b0;
            15'b11011100_1001_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 4 Row 10
            15'b11011100_1010_000: DATA = 1'b0;
            15'b11011100_1010_001: DATA = 1'b0;
            15'b11011100_1010_010: DATA = 1'b0;
            15'b11011100_1010_011: DATA = 1'b0;
            15'b11011100_1010_100: DATA = 1'b0;
            15'b11011100_1010_101: DATA = 1'b0;
            15'b11011100_1010_110: DATA = 1'b0;
            15'b11011100_1010_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 4 Row 11
            15'b11011100_1011_000: DATA = 1'b0;
            15'b11011100_1011_001: DATA = 1'b0;
            15'b11011100_1011_010: DATA = 1'b0;
            15'b11011100_1011_011: DATA = 1'b0;
            15'b11011100_1011_100: DATA = 1'b0;
            15'b11011100_1011_101: DATA = 1'b0;
            15'b11011100_1011_110: DATA = 1'b0;
            15'b11011100_1011_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 4 Row 12
            15'b11011100_1100_000: DATA = 1'b0;
            15'b11011100_1100_001: DATA = 1'b0;
            15'b11011100_1100_010: DATA = 1'b0;
            15'b11011100_1100_011: DATA = 1'b0;
            15'b11011100_1100_100: DATA = 1'b0;
            15'b11011100_1100_101: DATA = 1'b0;
            15'b11011100_1100_110: DATA = 1'b0;
            15'b11011100_1100_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 4 Row 13
            15'b11011100_1101_000: DATA = 1'b0;
            15'b11011100_1101_001: DATA = 1'b0;
            15'b11011100_1101_010: DATA = 1'b0;
            15'b11011100_1101_011: DATA = 1'b0;
            15'b11011100_1101_100: DATA = 1'b0;
            15'b11011100_1101_101: DATA = 1'b0;
            15'b11011100_1101_110: DATA = 1'b0;
            15'b11011100_1101_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 4 Row 14
            15'b11011100_1110_000: DATA = 1'b0;
            15'b11011100_1110_001: DATA = 1'b0;
            15'b11011100_1110_010: DATA = 1'b0;
            15'b11011100_1110_011: DATA = 1'b0;
            15'b11011100_1110_100: DATA = 1'b0;
            15'b11011100_1110_101: DATA = 1'b0;
            15'b11011100_1110_110: DATA = 1'b0;
            15'b11011100_1110_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 0 COL 4 Row 15
            15'b11011100_1111_000: DATA = 1'b0;
            15'b11011100_1111_001: DATA = 1'b0;
            15'b11011100_1111_010: DATA = 1'b0;
            15'b11011100_1111_011: DATA = 1'b0;
            15'b11011100_1111_100: DATA = 1'b0;
            15'b11011100_1111_101: DATA = 1'b0;
            15'b11011100_1111_110: DATA = 1'b0;
            15'b11011100_1111_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 0 Row 0
            15'b11011101_0000_000: DATA = 1'b1;
            15'b11011101_0000_001: DATA = 1'b0;
            15'b11011101_0000_010: DATA = 1'b0;
            15'b11011101_0000_011: DATA = 1'b0;
            15'b11011101_0000_100: DATA = 1'b0;
            15'b11011101_0000_101: DATA = 1'b0;
            15'b11011101_0000_110: DATA = 1'b0;
            15'b11011101_0000_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 0 Row 1
            15'b11011101_0001_000: DATA = 1'b1;
            15'b11011101_0001_001: DATA = 1'b0;
            15'b11011101_0001_010: DATA = 1'b0;
            15'b11011101_0001_011: DATA = 1'b0;
            15'b11011101_0001_100: DATA = 1'b0;
            15'b11011101_0001_101: DATA = 1'b0;
            15'b11011101_0001_110: DATA = 1'b0;
            15'b11011101_0001_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 0 Row 2
            15'b11011101_0010_000: DATA = 1'b1;
            15'b11011101_0010_001: DATA = 1'b0;
            15'b11011101_0010_010: DATA = 1'b0;
            15'b11011101_0010_011: DATA = 1'b0;
            15'b11011101_0010_100: DATA = 1'b0;
            15'b11011101_0010_101: DATA = 1'b0;
            15'b11011101_0010_110: DATA = 1'b0;
            15'b11011101_0010_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 0 Row 3
            15'b11011101_0011_000: DATA = 1'b1;
            15'b11011101_0011_001: DATA = 1'b0;
            15'b11011101_0011_010: DATA = 1'b0;
            15'b11011101_0011_011: DATA = 1'b0;
            15'b11011101_0011_100: DATA = 1'b0;
            15'b11011101_0011_101: DATA = 1'b0;
            15'b11011101_0011_110: DATA = 1'b0;
            15'b11011101_0011_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 0 Row 4
            15'b11011101_0100_000: DATA = 1'b1;
            15'b11011101_0100_001: DATA = 1'b0;
            15'b11011101_0100_010: DATA = 1'b0;
            15'b11011101_0100_011: DATA = 1'b0;
            15'b11011101_0100_100: DATA = 1'b0;
            15'b11011101_0100_101: DATA = 1'b0;
            15'b11011101_0100_110: DATA = 1'b0;
            15'b11011101_0100_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 0 Row 5
            15'b11011101_0101_000: DATA = 1'b1;
            15'b11011101_0101_001: DATA = 1'b0;
            15'b11011101_0101_010: DATA = 1'b0;
            15'b11011101_0101_011: DATA = 1'b0;
            15'b11011101_0101_100: DATA = 1'b0;
            15'b11011101_0101_101: DATA = 1'b0;
            15'b11011101_0101_110: DATA = 1'b0;
            15'b11011101_0101_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 0 Row 6
            15'b11011101_0110_000: DATA = 1'b1;
            15'b11011101_0110_001: DATA = 1'b0;
            15'b11011101_0110_010: DATA = 1'b0;
            15'b11011101_0110_011: DATA = 1'b0;
            15'b11011101_0110_100: DATA = 1'b0;
            15'b11011101_0110_101: DATA = 1'b0;
            15'b11011101_0110_110: DATA = 1'b0;
            15'b11011101_0110_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 0 Row 7
            15'b11011101_0111_000: DATA = 1'b1;
            15'b11011101_0111_001: DATA = 1'b0;
            15'b11011101_0111_010: DATA = 1'b0;
            15'b11011101_0111_011: DATA = 1'b0;
            15'b11011101_0111_100: DATA = 1'b0;
            15'b11011101_0111_101: DATA = 1'b0;
            15'b11011101_0111_110: DATA = 1'b0;
            15'b11011101_0111_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 0 Row 8
            15'b11011101_1000_000: DATA = 1'b1;
            15'b11011101_1000_001: DATA = 1'b0;
            15'b11011101_1000_010: DATA = 1'b0;
            15'b11011101_1000_011: DATA = 1'b0;
            15'b11011101_1000_100: DATA = 1'b0;
            15'b11011101_1000_101: DATA = 1'b0;
            15'b11011101_1000_110: DATA = 1'b0;
            15'b11011101_1000_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 0 Row 9
            15'b11011101_1001_000: DATA = 1'b1;
            15'b11011101_1001_001: DATA = 1'b0;
            15'b11011101_1001_010: DATA = 1'b0;
            15'b11011101_1001_011: DATA = 1'b0;
            15'b11011101_1001_100: DATA = 1'b0;
            15'b11011101_1001_101: DATA = 1'b0;
            15'b11011101_1001_110: DATA = 1'b0;
            15'b11011101_1001_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 0 Row 10
            15'b11011101_1010_000: DATA = 1'b1;
            15'b11011101_1010_001: DATA = 1'b0;
            15'b11011101_1010_010: DATA = 1'b0;
            15'b11011101_1010_011: DATA = 1'b0;
            15'b11011101_1010_100: DATA = 1'b0;
            15'b11011101_1010_101: DATA = 1'b0;
            15'b11011101_1010_110: DATA = 1'b0;
            15'b11011101_1010_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 0 Row 11
            15'b11011101_1011_000: DATA = 1'b1;
            15'b11011101_1011_001: DATA = 1'b0;
            15'b11011101_1011_010: DATA = 1'b0;
            15'b11011101_1011_011: DATA = 1'b0;
            15'b11011101_1011_100: DATA = 1'b0;
            15'b11011101_1011_101: DATA = 1'b0;
            15'b11011101_1011_110: DATA = 1'b0;
            15'b11011101_1011_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 0 Row 12
            15'b11011101_1100_000: DATA = 1'b1;
            15'b11011101_1100_001: DATA = 1'b0;
            15'b11011101_1100_010: DATA = 1'b0;
            15'b11011101_1100_011: DATA = 1'b0;
            15'b11011101_1100_100: DATA = 1'b0;
            15'b11011101_1100_101: DATA = 1'b0;
            15'b11011101_1100_110: DATA = 1'b0;
            15'b11011101_1100_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 0 Row 13
            15'b11011101_1101_000: DATA = 1'b1;
            15'b11011101_1101_001: DATA = 1'b0;
            15'b11011101_1101_010: DATA = 1'b0;
            15'b11011101_1101_011: DATA = 1'b0;
            15'b11011101_1101_100: DATA = 1'b0;
            15'b11011101_1101_101: DATA = 1'b0;
            15'b11011101_1101_110: DATA = 1'b0;
            15'b11011101_1101_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 0 Row 14
            15'b11011101_1110_000: DATA = 1'b1;
            15'b11011101_1110_001: DATA = 1'b0;
            15'b11011101_1110_010: DATA = 1'b0;
            15'b11011101_1110_011: DATA = 1'b0;
            15'b11011101_1110_100: DATA = 1'b0;
            15'b11011101_1110_101: DATA = 1'b0;
            15'b11011101_1110_110: DATA = 1'b0;
            15'b11011101_1110_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 0 Row 15
            15'b11011101_1111_000: DATA = 1'b1;
            15'b11011101_1111_001: DATA = 1'b0;
            15'b11011101_1111_010: DATA = 1'b0;
            15'b11011101_1111_011: DATA = 1'b0;
            15'b11011101_1111_100: DATA = 1'b0;
            15'b11011101_1111_101: DATA = 1'b0;
            15'b11011101_1111_110: DATA = 1'b0;
            15'b11011101_1111_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 1 Row 0
            15'b11011110_0000_000: DATA = 1'b0;
            15'b11011110_0000_001: DATA = 1'b0;
            15'b11011110_0000_010: DATA = 1'b0;
            15'b11011110_0000_011: DATA = 1'b0;
            15'b11011110_0000_100: DATA = 1'b0;
            15'b11011110_0000_101: DATA = 1'b0;
            15'b11011110_0000_110: DATA = 1'b0;
            15'b11011110_0000_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 1 Row 1
            15'b11011110_0001_000: DATA = 1'b0;
            15'b11011110_0001_001: DATA = 1'b0;
            15'b11011110_0001_010: DATA = 1'b0;
            15'b11011110_0001_011: DATA = 1'b0;
            15'b11011110_0001_100: DATA = 1'b0;
            15'b11011110_0001_101: DATA = 1'b0;
            15'b11011110_0001_110: DATA = 1'b0;
            15'b11011110_0001_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 1 Row 2
            15'b11011110_0010_000: DATA = 1'b0;
            15'b11011110_0010_001: DATA = 1'b0;
            15'b11011110_0010_010: DATA = 1'b0;
            15'b11011110_0010_011: DATA = 1'b0;
            15'b11011110_0010_100: DATA = 1'b0;
            15'b11011110_0010_101: DATA = 1'b0;
            15'b11011110_0010_110: DATA = 1'b0;
            15'b11011110_0010_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 1 Row 3
            15'b11011110_0011_000: DATA = 1'b0;
            15'b11011110_0011_001: DATA = 1'b0;
            15'b11011110_0011_010: DATA = 1'b0;
            15'b11011110_0011_011: DATA = 1'b0;
            15'b11011110_0011_100: DATA = 1'b0;
            15'b11011110_0011_101: DATA = 1'b0;
            15'b11011110_0011_110: DATA = 1'b0;
            15'b11011110_0011_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 1 Row 4
            15'b11011110_0100_000: DATA = 1'b0;
            15'b11011110_0100_001: DATA = 1'b0;
            15'b11011110_0100_010: DATA = 1'b0;
            15'b11011110_0100_011: DATA = 1'b0;
            15'b11011110_0100_100: DATA = 1'b0;
            15'b11011110_0100_101: DATA = 1'b0;
            15'b11011110_0100_110: DATA = 1'b0;
            15'b11011110_0100_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 1 Row 5
            15'b11011110_0101_000: DATA = 1'b0;
            15'b11011110_0101_001: DATA = 1'b0;
            15'b11011110_0101_010: DATA = 1'b0;
            15'b11011110_0101_011: DATA = 1'b0;
            15'b11011110_0101_100: DATA = 1'b0;
            15'b11011110_0101_101: DATA = 1'b0;
            15'b11011110_0101_110: DATA = 1'b0;
            15'b11011110_0101_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 1 Row 6
            15'b11011110_0110_000: DATA = 1'b0;
            15'b11011110_0110_001: DATA = 1'b0;
            15'b11011110_0110_010: DATA = 1'b0;
            15'b11011110_0110_011: DATA = 1'b0;
            15'b11011110_0110_100: DATA = 1'b0;
            15'b11011110_0110_101: DATA = 1'b0;
            15'b11011110_0110_110: DATA = 1'b0;
            15'b11011110_0110_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 1 Row 7
            15'b11011110_0111_000: DATA = 1'b0;
            15'b11011110_0111_001: DATA = 1'b0;
            15'b11011110_0111_010: DATA = 1'b0;
            15'b11011110_0111_011: DATA = 1'b0;
            15'b11011110_0111_100: DATA = 1'b0;
            15'b11011110_0111_101: DATA = 1'b0;
            15'b11011110_0111_110: DATA = 1'b0;
            15'b11011110_0111_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 1 Row 8
            15'b11011110_1000_000: DATA = 1'b0;
            15'b11011110_1000_001: DATA = 1'b0;
            15'b11011110_1000_010: DATA = 1'b0;
            15'b11011110_1000_011: DATA = 1'b0;
            15'b11011110_1000_100: DATA = 1'b0;
            15'b11011110_1000_101: DATA = 1'b0;
            15'b11011110_1000_110: DATA = 1'b0;
            15'b11011110_1000_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 1 Row 9
            15'b11011110_1001_000: DATA = 1'b0;
            15'b11011110_1001_001: DATA = 1'b0;
            15'b11011110_1001_010: DATA = 1'b0;
            15'b11011110_1001_011: DATA = 1'b0;
            15'b11011110_1001_100: DATA = 1'b0;
            15'b11011110_1001_101: DATA = 1'b0;
            15'b11011110_1001_110: DATA = 1'b0;
            15'b11011110_1001_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 1 Row 10
            15'b11011110_1010_000: DATA = 1'b0;
            15'b11011110_1010_001: DATA = 1'b0;
            15'b11011110_1010_010: DATA = 1'b0;
            15'b11011110_1010_011: DATA = 1'b0;
            15'b11011110_1010_100: DATA = 1'b0;
            15'b11011110_1010_101: DATA = 1'b0;
            15'b11011110_1010_110: DATA = 1'b0;
            15'b11011110_1010_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 1 Row 11
            15'b11011110_1011_000: DATA = 1'b0;
            15'b11011110_1011_001: DATA = 1'b0;
            15'b11011110_1011_010: DATA = 1'b0;
            15'b11011110_1011_011: DATA = 1'b0;
            15'b11011110_1011_100: DATA = 1'b0;
            15'b11011110_1011_101: DATA = 1'b0;
            15'b11011110_1011_110: DATA = 1'b0;
            15'b11011110_1011_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 1 Row 12
            15'b11011110_1100_000: DATA = 1'b0;
            15'b11011110_1100_001: DATA = 1'b0;
            15'b11011110_1100_010: DATA = 1'b0;
            15'b11011110_1100_011: DATA = 1'b0;
            15'b11011110_1100_100: DATA = 1'b0;
            15'b11011110_1100_101: DATA = 1'b0;
            15'b11011110_1100_110: DATA = 1'b0;
            15'b11011110_1100_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 1 Row 13
            15'b11011110_1101_000: DATA = 1'b0;
            15'b11011110_1101_001: DATA = 1'b0;
            15'b11011110_1101_010: DATA = 1'b0;
            15'b11011110_1101_011: DATA = 1'b0;
            15'b11011110_1101_100: DATA = 1'b0;
            15'b11011110_1101_101: DATA = 1'b0;
            15'b11011110_1101_110: DATA = 1'b0;
            15'b11011110_1101_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 1 Row 14
            15'b11011110_1110_000: DATA = 1'b0;
            15'b11011110_1110_001: DATA = 1'b0;
            15'b11011110_1110_010: DATA = 1'b0;
            15'b11011110_1110_011: DATA = 1'b0;
            15'b11011110_1110_100: DATA = 1'b0;
            15'b11011110_1110_101: DATA = 1'b0;
            15'b11011110_1110_110: DATA = 1'b0;
            15'b11011110_1110_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 1 Row 15
            15'b11011110_1111_000: DATA = 1'b0;
            15'b11011110_1111_001: DATA = 1'b0;
            15'b11011110_1111_010: DATA = 1'b0;
            15'b11011110_1111_011: DATA = 1'b0;
            15'b11011110_1111_100: DATA = 1'b0;
            15'b11011110_1111_101: DATA = 1'b0;
            15'b11011110_1111_110: DATA = 1'b0;
            15'b11011110_1111_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 2 Row 0
            15'b11011111_0000_000: DATA = 1'b0;
            15'b11011111_0000_001: DATA = 1'b0;
            15'b11011111_0000_010: DATA = 1'b0;
            15'b11011111_0000_011: DATA = 1'b1;
            15'b11011111_0000_100: DATA = 1'b1;
            15'b11011111_0000_101: DATA = 1'b1;
            15'b11011111_0000_110: DATA = 1'b0;
            15'b11011111_0000_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 2 Row 1
            15'b11011111_0001_000: DATA = 1'b0;
            15'b11011111_0001_001: DATA = 1'b0;
            15'b11011111_0001_010: DATA = 1'b0;
            15'b11011111_0001_011: DATA = 1'b0;
            15'b11011111_0001_100: DATA = 1'b0;
            15'b11011111_0001_101: DATA = 1'b1;
            15'b11011111_0001_110: DATA = 1'b1;
            15'b11011111_0001_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 2 Row 2
            15'b11011111_0010_000: DATA = 1'b0;
            15'b11011111_0010_001: DATA = 1'b0;
            15'b11011111_0010_010: DATA = 1'b0;
            15'b11011111_0010_011: DATA = 1'b0;
            15'b11011111_0010_100: DATA = 1'b0;
            15'b11011111_0010_101: DATA = 1'b0;
            15'b11011111_0010_110: DATA = 1'b1;
            15'b11011111_0010_111: DATA = 1'b1;
            //SAWTOOTHY+ ROW 1 COL 2 Row 3
            15'b11011111_0011_000: DATA = 1'b0;
            15'b11011111_0011_001: DATA = 1'b0;
            15'b11011111_0011_010: DATA = 1'b0;
            15'b11011111_0011_011: DATA = 1'b0;
            15'b11011111_0011_100: DATA = 1'b0;
            15'b11011111_0011_101: DATA = 1'b0;
            15'b11011111_0011_110: DATA = 1'b0;
            15'b11011111_0011_111: DATA = 1'b1;
            //SAWTOOTHY+ ROW 1 COL 2 Row 4
            15'b11011111_0100_000: DATA = 1'b0;
            15'b11011111_0100_001: DATA = 1'b0;
            15'b11011111_0100_010: DATA = 1'b0;
            15'b11011111_0100_011: DATA = 1'b0;
            15'b11011111_0100_100: DATA = 1'b0;
            15'b11011111_0100_101: DATA = 1'b0;
            15'b11011111_0100_110: DATA = 1'b0;
            15'b11011111_0100_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 2 Row 5
            15'b11011111_0101_000: DATA = 1'b0;
            15'b11011111_0101_001: DATA = 1'b0;
            15'b11011111_0101_010: DATA = 1'b0;
            15'b11011111_0101_011: DATA = 1'b0;
            15'b11011111_0101_100: DATA = 1'b0;
            15'b11011111_0101_101: DATA = 1'b0;
            15'b11011111_0101_110: DATA = 1'b0;
            15'b11011111_0101_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 2 Row 6
            15'b11011111_0110_000: DATA = 1'b0;
            15'b11011111_0110_001: DATA = 1'b0;
            15'b11011111_0110_010: DATA = 1'b0;
            15'b11011111_0110_011: DATA = 1'b0;
            15'b11011111_0110_100: DATA = 1'b0;
            15'b11011111_0110_101: DATA = 1'b0;
            15'b11011111_0110_110: DATA = 1'b0;
            15'b11011111_0110_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 2 Row 7
            15'b11011111_0111_000: DATA = 1'b0;
            15'b11011111_0111_001: DATA = 1'b0;
            15'b11011111_0111_010: DATA = 1'b0;
            15'b11011111_0111_011: DATA = 1'b0;
            15'b11011111_0111_100: DATA = 1'b0;
            15'b11011111_0111_101: DATA = 1'b0;
            15'b11011111_0111_110: DATA = 1'b0;
            15'b11011111_0111_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 2 Row 8
            15'b11011111_1000_000: DATA = 1'b0;
            15'b11011111_1000_001: DATA = 1'b0;
            15'b11011111_1000_010: DATA = 1'b0;
            15'b11011111_1000_011: DATA = 1'b0;
            15'b11011111_1000_100: DATA = 1'b0;
            15'b11011111_1000_101: DATA = 1'b0;
            15'b11011111_1000_110: DATA = 1'b0;
            15'b11011111_1000_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 2 Row 9
            15'b11011111_1001_000: DATA = 1'b0;
            15'b11011111_1001_001: DATA = 1'b0;
            15'b11011111_1001_010: DATA = 1'b0;
            15'b11011111_1001_011: DATA = 1'b0;
            15'b11011111_1001_100: DATA = 1'b0;
            15'b11011111_1001_101: DATA = 1'b0;
            15'b11011111_1001_110: DATA = 1'b0;
            15'b11011111_1001_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 2 Row 10
            15'b11011111_1010_000: DATA = 1'b0;
            15'b11011111_1010_001: DATA = 1'b0;
            15'b11011111_1010_010: DATA = 1'b0;
            15'b11011111_1010_011: DATA = 1'b0;
            15'b11011111_1010_100: DATA = 1'b0;
            15'b11011111_1010_101: DATA = 1'b0;
            15'b11011111_1010_110: DATA = 1'b0;
            15'b11011111_1010_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 2 Row 11
            15'b11011111_1011_000: DATA = 1'b0;
            15'b11011111_1011_001: DATA = 1'b0;
            15'b11011111_1011_010: DATA = 1'b0;
            15'b11011111_1011_011: DATA = 1'b0;
            15'b11011111_1011_100: DATA = 1'b0;
            15'b11011111_1011_101: DATA = 1'b0;
            15'b11011111_1011_110: DATA = 1'b0;
            15'b11011111_1011_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 2 Row 12
            15'b11011111_1100_000: DATA = 1'b0;
            15'b11011111_1100_001: DATA = 1'b0;
            15'b11011111_1100_010: DATA = 1'b0;
            15'b11011111_1100_011: DATA = 1'b0;
            15'b11011111_1100_100: DATA = 1'b0;
            15'b11011111_1100_101: DATA = 1'b0;
            15'b11011111_1100_110: DATA = 1'b0;
            15'b11011111_1100_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 2 Row 13
            15'b11011111_1101_000: DATA = 1'b0;
            15'b11011111_1101_001: DATA = 1'b0;
            15'b11011111_1101_010: DATA = 1'b0;
            15'b11011111_1101_011: DATA = 1'b0;
            15'b11011111_1101_100: DATA = 1'b0;
            15'b11011111_1101_101: DATA = 1'b0;
            15'b11011111_1101_110: DATA = 1'b0;
            15'b11011111_1101_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 2 Row 14
            15'b11011111_1110_000: DATA = 1'b0;
            15'b11011111_1110_001: DATA = 1'b0;
            15'b11011111_1110_010: DATA = 1'b0;
            15'b11011111_1110_011: DATA = 1'b0;
            15'b11011111_1110_100: DATA = 1'b0;
            15'b11011111_1110_101: DATA = 1'b0;
            15'b11011111_1110_110: DATA = 1'b0;
            15'b11011111_1110_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 2 Row 15
            15'b11011111_1111_000: DATA = 1'b0;
            15'b11011111_1111_001: DATA = 1'b0;
            15'b11011111_1111_010: DATA = 1'b0;
            15'b11011111_1111_011: DATA = 1'b0;
            15'b11011111_1111_100: DATA = 1'b0;
            15'b11011111_1111_101: DATA = 1'b0;
            15'b11011111_1111_110: DATA = 1'b0;
            15'b11011111_1111_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 3 Row 0
            15'b11100000_0000_000: DATA = 1'b0;
            15'b11100000_0000_001: DATA = 1'b0;
            15'b11100000_0000_010: DATA = 1'b0;
            15'b11100000_0000_011: DATA = 1'b0;
            15'b11100000_0000_100: DATA = 1'b0;
            15'b11100000_0000_101: DATA = 1'b0;
            15'b11100000_0000_110: DATA = 1'b0;
            15'b11100000_0000_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 3 Row 1
            15'b11100000_0001_000: DATA = 1'b0;
            15'b11100000_0001_001: DATA = 1'b0;
            15'b11100000_0001_010: DATA = 1'b0;
            15'b11100000_0001_011: DATA = 1'b0;
            15'b11100000_0001_100: DATA = 1'b0;
            15'b11100000_0001_101: DATA = 1'b0;
            15'b11100000_0001_110: DATA = 1'b0;
            15'b11100000_0001_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 3 Row 2
            15'b11100000_0010_000: DATA = 1'b0;
            15'b11100000_0010_001: DATA = 1'b0;
            15'b11100000_0010_010: DATA = 1'b0;
            15'b11100000_0010_011: DATA = 1'b0;
            15'b11100000_0010_100: DATA = 1'b0;
            15'b11100000_0010_101: DATA = 1'b0;
            15'b11100000_0010_110: DATA = 1'b0;
            15'b11100000_0010_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 3 Row 3
            15'b11100000_0011_000: DATA = 1'b1;
            15'b11100000_0011_001: DATA = 1'b0;
            15'b11100000_0011_010: DATA = 1'b0;
            15'b11100000_0011_011: DATA = 1'b0;
            15'b11100000_0011_100: DATA = 1'b0;
            15'b11100000_0011_101: DATA = 1'b0;
            15'b11100000_0011_110: DATA = 1'b0;
            15'b11100000_0011_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 3 Row 4
            15'b11100000_0100_000: DATA = 1'b1;
            15'b11100000_0100_001: DATA = 1'b1;
            15'b11100000_0100_010: DATA = 1'b1;
            15'b11100000_0100_011: DATA = 1'b0;
            15'b11100000_0100_100: DATA = 1'b0;
            15'b11100000_0100_101: DATA = 1'b0;
            15'b11100000_0100_110: DATA = 1'b0;
            15'b11100000_0100_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 3 Row 5
            15'b11100000_0101_000: DATA = 1'b0;
            15'b11100000_0101_001: DATA = 1'b0;
            15'b11100000_0101_010: DATA = 1'b1;
            15'b11100000_0101_011: DATA = 1'b1;
            15'b11100000_0101_100: DATA = 1'b0;
            15'b11100000_0101_101: DATA = 1'b0;
            15'b11100000_0101_110: DATA = 1'b0;
            15'b11100000_0101_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 3 Row 6
            15'b11100000_0110_000: DATA = 1'b0;
            15'b11100000_0110_001: DATA = 1'b0;
            15'b11100000_0110_010: DATA = 1'b0;
            15'b11100000_0110_011: DATA = 1'b1;
            15'b11100000_0110_100: DATA = 1'b1;
            15'b11100000_0110_101: DATA = 1'b0;
            15'b11100000_0110_110: DATA = 1'b0;
            15'b11100000_0110_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 3 Row 7
            15'b11100000_0111_000: DATA = 1'b0;
            15'b11100000_0111_001: DATA = 1'b0;
            15'b11100000_0111_010: DATA = 1'b0;
            15'b11100000_0111_011: DATA = 1'b0;
            15'b11100000_0111_100: DATA = 1'b1;
            15'b11100000_0111_101: DATA = 1'b1;
            15'b11100000_0111_110: DATA = 1'b0;
            15'b11100000_0111_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 3 Row 8
            15'b11100000_1000_000: DATA = 1'b0;
            15'b11100000_1000_001: DATA = 1'b0;
            15'b11100000_1000_010: DATA = 1'b0;
            15'b11100000_1000_011: DATA = 1'b0;
            15'b11100000_1000_100: DATA = 1'b0;
            15'b11100000_1000_101: DATA = 1'b1;
            15'b11100000_1000_110: DATA = 1'b1;
            15'b11100000_1000_111: DATA = 1'b1;
            //SAWTOOTHY+ ROW 1 COL 3 Row 9
            15'b11100000_1001_000: DATA = 1'b0;
            15'b11100000_1001_001: DATA = 1'b0;
            15'b11100000_1001_010: DATA = 1'b0;
            15'b11100000_1001_011: DATA = 1'b0;
            15'b11100000_1001_100: DATA = 1'b0;
            15'b11100000_1001_101: DATA = 1'b0;
            15'b11100000_1001_110: DATA = 1'b0;
            15'b11100000_1001_111: DATA = 1'b1;
            //SAWTOOTHY+ ROW 1 COL 3 Row 10
            15'b11100000_1010_000: DATA = 1'b0;
            15'b11100000_1010_001: DATA = 1'b0;
            15'b11100000_1010_010: DATA = 1'b0;
            15'b11100000_1010_011: DATA = 1'b0;
            15'b11100000_1010_100: DATA = 1'b0;
            15'b11100000_1010_101: DATA = 1'b0;
            15'b11100000_1010_110: DATA = 1'b0;
            15'b11100000_1010_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 3 Row 11
            15'b11100000_1011_000: DATA = 1'b0;
            15'b11100000_1011_001: DATA = 1'b0;
            15'b11100000_1011_010: DATA = 1'b0;
            15'b11100000_1011_011: DATA = 1'b0;
            15'b11100000_1011_100: DATA = 1'b0;
            15'b11100000_1011_101: DATA = 1'b0;
            15'b11100000_1011_110: DATA = 1'b0;
            15'b11100000_1011_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 3 Row 12
            15'b11100000_1100_000: DATA = 1'b0;
            15'b11100000_1100_001: DATA = 1'b0;
            15'b11100000_1100_010: DATA = 1'b0;
            15'b11100000_1100_011: DATA = 1'b0;
            15'b11100000_1100_100: DATA = 1'b0;
            15'b11100000_1100_101: DATA = 1'b0;
            15'b11100000_1100_110: DATA = 1'b0;
            15'b11100000_1100_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 3 Row 13
            15'b11100000_1101_000: DATA = 1'b0;
            15'b11100000_1101_001: DATA = 1'b0;
            15'b11100000_1101_010: DATA = 1'b0;
            15'b11100000_1101_011: DATA = 1'b0;
            15'b11100000_1101_100: DATA = 1'b0;
            15'b11100000_1101_101: DATA = 1'b0;
            15'b11100000_1101_110: DATA = 1'b0;
            15'b11100000_1101_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 3 Row 14
            15'b11100000_1110_000: DATA = 1'b0;
            15'b11100000_1110_001: DATA = 1'b0;
            15'b11100000_1110_010: DATA = 1'b0;
            15'b11100000_1110_011: DATA = 1'b0;
            15'b11100000_1110_100: DATA = 1'b0;
            15'b11100000_1110_101: DATA = 1'b0;
            15'b11100000_1110_110: DATA = 1'b0;
            15'b11100000_1110_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 3 Row 15
            15'b11100000_1111_000: DATA = 1'b0;
            15'b11100000_1111_001: DATA = 1'b0;
            15'b11100000_1111_010: DATA = 1'b0;
            15'b11100000_1111_011: DATA = 1'b0;
            15'b11100000_1111_100: DATA = 1'b0;
            15'b11100000_1111_101: DATA = 1'b0;
            15'b11100000_1111_110: DATA = 1'b0;
            15'b11100000_1111_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 4 Row 0
            15'b11100001_0000_000: DATA = 1'b0;
            15'b11100001_0000_001: DATA = 1'b0;
            15'b11100001_0000_010: DATA = 1'b0;
            15'b11100001_0000_011: DATA = 1'b0;
            15'b11100001_0000_100: DATA = 1'b0;
            15'b11100001_0000_101: DATA = 1'b0;
            15'b11100001_0000_110: DATA = 1'b0;
            15'b11100001_0000_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 4 Row 1
            15'b11100001_0001_000: DATA = 1'b0;
            15'b11100001_0001_001: DATA = 1'b0;
            15'b11100001_0001_010: DATA = 1'b0;
            15'b11100001_0001_011: DATA = 1'b0;
            15'b11100001_0001_100: DATA = 1'b0;
            15'b11100001_0001_101: DATA = 1'b0;
            15'b11100001_0001_110: DATA = 1'b0;
            15'b11100001_0001_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 4 Row 2
            15'b11100001_0010_000: DATA = 1'b0;
            15'b11100001_0010_001: DATA = 1'b0;
            15'b11100001_0010_010: DATA = 1'b0;
            15'b11100001_0010_011: DATA = 1'b0;
            15'b11100001_0010_100: DATA = 1'b0;
            15'b11100001_0010_101: DATA = 1'b0;
            15'b11100001_0010_110: DATA = 1'b0;
            15'b11100001_0010_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 4 Row 3
            15'b11100001_0011_000: DATA = 1'b0;
            15'b11100001_0011_001: DATA = 1'b0;
            15'b11100001_0011_010: DATA = 1'b0;
            15'b11100001_0011_011: DATA = 1'b0;
            15'b11100001_0011_100: DATA = 1'b0;
            15'b11100001_0011_101: DATA = 1'b0;
            15'b11100001_0011_110: DATA = 1'b0;
            15'b11100001_0011_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 4 Row 4
            15'b11100001_0100_000: DATA = 1'b0;
            15'b11100001_0100_001: DATA = 1'b0;
            15'b11100001_0100_010: DATA = 1'b0;
            15'b11100001_0100_011: DATA = 1'b0;
            15'b11100001_0100_100: DATA = 1'b0;
            15'b11100001_0100_101: DATA = 1'b0;
            15'b11100001_0100_110: DATA = 1'b0;
            15'b11100001_0100_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 4 Row 5
            15'b11100001_0101_000: DATA = 1'b0;
            15'b11100001_0101_001: DATA = 1'b0;
            15'b11100001_0101_010: DATA = 1'b0;
            15'b11100001_0101_011: DATA = 1'b0;
            15'b11100001_0101_100: DATA = 1'b0;
            15'b11100001_0101_101: DATA = 1'b0;
            15'b11100001_0101_110: DATA = 1'b0;
            15'b11100001_0101_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 4 Row 6
            15'b11100001_0110_000: DATA = 1'b0;
            15'b11100001_0110_001: DATA = 1'b0;
            15'b11100001_0110_010: DATA = 1'b0;
            15'b11100001_0110_011: DATA = 1'b0;
            15'b11100001_0110_100: DATA = 1'b0;
            15'b11100001_0110_101: DATA = 1'b0;
            15'b11100001_0110_110: DATA = 1'b0;
            15'b11100001_0110_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 4 Row 7
            15'b11100001_0111_000: DATA = 1'b0;
            15'b11100001_0111_001: DATA = 1'b0;
            15'b11100001_0111_010: DATA = 1'b0;
            15'b11100001_0111_011: DATA = 1'b0;
            15'b11100001_0111_100: DATA = 1'b0;
            15'b11100001_0111_101: DATA = 1'b0;
            15'b11100001_0111_110: DATA = 1'b0;
            15'b11100001_0111_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 4 Row 8
            15'b11100001_1000_000: DATA = 1'b0;
            15'b11100001_1000_001: DATA = 1'b0;
            15'b11100001_1000_010: DATA = 1'b0;
            15'b11100001_1000_011: DATA = 1'b0;
            15'b11100001_1000_100: DATA = 1'b0;
            15'b11100001_1000_101: DATA = 1'b0;
            15'b11100001_1000_110: DATA = 1'b0;
            15'b11100001_1000_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 4 Row 9
            15'b11100001_1001_000: DATA = 1'b1;
            15'b11100001_1001_001: DATA = 1'b0;
            15'b11100001_1001_010: DATA = 1'b0;
            15'b11100001_1001_011: DATA = 1'b0;
            15'b11100001_1001_100: DATA = 1'b0;
            15'b11100001_1001_101: DATA = 1'b0;
            15'b11100001_1001_110: DATA = 1'b0;
            15'b11100001_1001_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 4 Row 10
            15'b11100001_1010_000: DATA = 1'b1;
            15'b11100001_1010_001: DATA = 1'b1;
            15'b11100001_1010_010: DATA = 1'b0;
            15'b11100001_1010_011: DATA = 1'b0;
            15'b11100001_1010_100: DATA = 1'b0;
            15'b11100001_1010_101: DATA = 1'b0;
            15'b11100001_1010_110: DATA = 1'b0;
            15'b11100001_1010_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 4 Row 11
            15'b11100001_1011_000: DATA = 1'b0;
            15'b11100001_1011_001: DATA = 1'b1;
            15'b11100001_1011_010: DATA = 1'b1;
            15'b11100001_1011_011: DATA = 1'b0;
            15'b11100001_1011_100: DATA = 1'b0;
            15'b11100001_1011_101: DATA = 1'b0;
            15'b11100001_1011_110: DATA = 1'b0;
            15'b11100001_1011_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 4 Row 12
            15'b11100001_1100_000: DATA = 1'b0;
            15'b11100001_1100_001: DATA = 1'b0;
            15'b11100001_1100_010: DATA = 1'b1;
            15'b11100001_1100_011: DATA = 1'b1;
            15'b11100001_1100_100: DATA = 1'b1;
            15'b11100001_1100_101: DATA = 1'b0;
            15'b11100001_1100_110: DATA = 1'b0;
            15'b11100001_1100_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 4 Row 13
            15'b11100001_1101_000: DATA = 1'b0;
            15'b11100001_1101_001: DATA = 1'b0;
            15'b11100001_1101_010: DATA = 1'b0;
            15'b11100001_1101_011: DATA = 1'b0;
            15'b11100001_1101_100: DATA = 1'b1;
            15'b11100001_1101_101: DATA = 1'b1;
            15'b11100001_1101_110: DATA = 1'b0;
            15'b11100001_1101_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 4 Row 14
            15'b11100001_1110_000: DATA = 1'b0;
            15'b11100001_1110_001: DATA = 1'b0;
            15'b11100001_1110_010: DATA = 1'b0;
            15'b11100001_1110_011: DATA = 1'b0;
            15'b11100001_1110_100: DATA = 1'b0;
            15'b11100001_1110_101: DATA = 1'b1;
            15'b11100001_1110_110: DATA = 1'b1;
            15'b11100001_1110_111: DATA = 1'b0;
            //SAWTOOTHY+ ROW 1 COL 4 Row 15
            15'b11100001_1111_000: DATA = 1'b0;
            15'b11100001_1111_001: DATA = 1'b0;
            15'b11100001_1111_010: DATA = 1'b0;
            15'b11100001_1111_011: DATA = 1'b0;
            15'b11100001_1111_100: DATA = 1'b0;
            15'b11100001_1111_101: DATA = 1'b0;
            15'b11100001_1111_110: DATA = 1'b1;
            15'b11100001_1111_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 0 COL 0 Row 0
            15'b11100010_0000_000: DATA = 1'b1;
            15'b11100010_0000_001: DATA = 1'b1;
            15'b11100010_0000_010: DATA = 1'b0;
            15'b11100010_0000_011: DATA = 1'b0;
            15'b11100010_0000_100: DATA = 1'b0;
            15'b11100010_0000_101: DATA = 1'b0;
            15'b11100010_0000_110: DATA = 1'b0;
            15'b11100010_0000_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 0 Row 1
            15'b11100010_0001_000: DATA = 1'b0;
            15'b11100010_0001_001: DATA = 1'b1;
            15'b11100010_0001_010: DATA = 1'b1;
            15'b11100010_0001_011: DATA = 1'b0;
            15'b11100010_0001_100: DATA = 1'b0;
            15'b11100010_0001_101: DATA = 1'b0;
            15'b11100010_0001_110: DATA = 1'b0;
            15'b11100010_0001_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 0 Row 2
            15'b11100010_0010_000: DATA = 1'b0;
            15'b11100010_0010_001: DATA = 1'b0;
            15'b11100010_0010_010: DATA = 1'b1;
            15'b11100010_0010_011: DATA = 1'b1;
            15'b11100010_0010_100: DATA = 1'b0;
            15'b11100010_0010_101: DATA = 1'b0;
            15'b11100010_0010_110: DATA = 1'b0;
            15'b11100010_0010_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 0 Row 3
            15'b11100010_0011_000: DATA = 1'b0;
            15'b11100010_0011_001: DATA = 1'b0;
            15'b11100010_0011_010: DATA = 1'b0;
            15'b11100010_0011_011: DATA = 1'b1;
            15'b11100010_0011_100: DATA = 1'b1;
            15'b11100010_0011_101: DATA = 1'b1;
            15'b11100010_0011_110: DATA = 1'b0;
            15'b11100010_0011_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 0 Row 4
            15'b11100010_0100_000: DATA = 1'b0;
            15'b11100010_0100_001: DATA = 1'b0;
            15'b11100010_0100_010: DATA = 1'b0;
            15'b11100010_0100_011: DATA = 1'b0;
            15'b11100010_0100_100: DATA = 1'b0;
            15'b11100010_0100_101: DATA = 1'b1;
            15'b11100010_0100_110: DATA = 1'b1;
            15'b11100010_0100_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 0 Row 5
            15'b11100010_0101_000: DATA = 1'b0;
            15'b11100010_0101_001: DATA = 1'b0;
            15'b11100010_0101_010: DATA = 1'b0;
            15'b11100010_0101_011: DATA = 1'b0;
            15'b11100010_0101_100: DATA = 1'b0;
            15'b11100010_0101_101: DATA = 1'b0;
            15'b11100010_0101_110: DATA = 1'b1;
            15'b11100010_0101_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 0 COL 0 Row 6
            15'b11100010_0110_000: DATA = 1'b0;
            15'b11100010_0110_001: DATA = 1'b0;
            15'b11100010_0110_010: DATA = 1'b0;
            15'b11100010_0110_011: DATA = 1'b0;
            15'b11100010_0110_100: DATA = 1'b0;
            15'b11100010_0110_101: DATA = 1'b0;
            15'b11100010_0110_110: DATA = 1'b0;
            15'b11100010_0110_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 0 COL 0 Row 7
            15'b11100010_0111_000: DATA = 1'b0;
            15'b11100010_0111_001: DATA = 1'b0;
            15'b11100010_0111_010: DATA = 1'b0;
            15'b11100010_0111_011: DATA = 1'b0;
            15'b11100010_0111_100: DATA = 1'b0;
            15'b11100010_0111_101: DATA = 1'b0;
            15'b11100010_0111_110: DATA = 1'b0;
            15'b11100010_0111_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 0 Row 8
            15'b11100010_1000_000: DATA = 1'b0;
            15'b11100010_1000_001: DATA = 1'b0;
            15'b11100010_1000_010: DATA = 1'b0;
            15'b11100010_1000_011: DATA = 1'b0;
            15'b11100010_1000_100: DATA = 1'b0;
            15'b11100010_1000_101: DATA = 1'b0;
            15'b11100010_1000_110: DATA = 1'b0;
            15'b11100010_1000_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 0 Row 9
            15'b11100010_1001_000: DATA = 1'b0;
            15'b11100010_1001_001: DATA = 1'b0;
            15'b11100010_1001_010: DATA = 1'b0;
            15'b11100010_1001_011: DATA = 1'b0;
            15'b11100010_1001_100: DATA = 1'b0;
            15'b11100010_1001_101: DATA = 1'b0;
            15'b11100010_1001_110: DATA = 1'b0;
            15'b11100010_1001_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 0 Row 10
            15'b11100010_1010_000: DATA = 1'b0;
            15'b11100010_1010_001: DATA = 1'b0;
            15'b11100010_1010_010: DATA = 1'b0;
            15'b11100010_1010_011: DATA = 1'b0;
            15'b11100010_1010_100: DATA = 1'b0;
            15'b11100010_1010_101: DATA = 1'b0;
            15'b11100010_1010_110: DATA = 1'b0;
            15'b11100010_1010_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 0 Row 11
            15'b11100010_1011_000: DATA = 1'b0;
            15'b11100010_1011_001: DATA = 1'b0;
            15'b11100010_1011_010: DATA = 1'b0;
            15'b11100010_1011_011: DATA = 1'b0;
            15'b11100010_1011_100: DATA = 1'b0;
            15'b11100010_1011_101: DATA = 1'b0;
            15'b11100010_1011_110: DATA = 1'b0;
            15'b11100010_1011_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 0 Row 12
            15'b11100010_1100_000: DATA = 1'b0;
            15'b11100010_1100_001: DATA = 1'b0;
            15'b11100010_1100_010: DATA = 1'b0;
            15'b11100010_1100_011: DATA = 1'b0;
            15'b11100010_1100_100: DATA = 1'b0;
            15'b11100010_1100_101: DATA = 1'b0;
            15'b11100010_1100_110: DATA = 1'b0;
            15'b11100010_1100_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 0 Row 13
            15'b11100010_1101_000: DATA = 1'b0;
            15'b11100010_1101_001: DATA = 1'b0;
            15'b11100010_1101_010: DATA = 1'b0;
            15'b11100010_1101_011: DATA = 1'b0;
            15'b11100010_1101_100: DATA = 1'b0;
            15'b11100010_1101_101: DATA = 1'b0;
            15'b11100010_1101_110: DATA = 1'b0;
            15'b11100010_1101_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 0 Row 14
            15'b11100010_1110_000: DATA = 1'b0;
            15'b11100010_1110_001: DATA = 1'b0;
            15'b11100010_1110_010: DATA = 1'b0;
            15'b11100010_1110_011: DATA = 1'b0;
            15'b11100010_1110_100: DATA = 1'b0;
            15'b11100010_1110_101: DATA = 1'b0;
            15'b11100010_1110_110: DATA = 1'b0;
            15'b11100010_1110_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 0 Row 15
            15'b11100010_1111_000: DATA = 1'b0;
            15'b11100010_1111_001: DATA = 1'b0;
            15'b11100010_1111_010: DATA = 1'b0;
            15'b11100010_1111_011: DATA = 1'b0;
            15'b11100010_1111_100: DATA = 1'b0;
            15'b11100010_1111_101: DATA = 1'b0;
            15'b11100010_1111_110: DATA = 1'b0;
            15'b11100010_1111_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 1 Row 0
            15'b11100011_0000_000: DATA = 1'b0;
            15'b11100011_0000_001: DATA = 1'b0;
            15'b11100011_0000_010: DATA = 1'b0;
            15'b11100011_0000_011: DATA = 1'b0;
            15'b11100011_0000_100: DATA = 1'b0;
            15'b11100011_0000_101: DATA = 1'b0;
            15'b11100011_0000_110: DATA = 1'b0;
            15'b11100011_0000_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 1 Row 1
            15'b11100011_0001_000: DATA = 1'b0;
            15'b11100011_0001_001: DATA = 1'b0;
            15'b11100011_0001_010: DATA = 1'b0;
            15'b11100011_0001_011: DATA = 1'b0;
            15'b11100011_0001_100: DATA = 1'b0;
            15'b11100011_0001_101: DATA = 1'b0;
            15'b11100011_0001_110: DATA = 1'b0;
            15'b11100011_0001_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 1 Row 2
            15'b11100011_0010_000: DATA = 1'b0;
            15'b11100011_0010_001: DATA = 1'b0;
            15'b11100011_0010_010: DATA = 1'b0;
            15'b11100011_0010_011: DATA = 1'b0;
            15'b11100011_0010_100: DATA = 1'b0;
            15'b11100011_0010_101: DATA = 1'b0;
            15'b11100011_0010_110: DATA = 1'b0;
            15'b11100011_0010_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 1 Row 3
            15'b11100011_0011_000: DATA = 1'b0;
            15'b11100011_0011_001: DATA = 1'b0;
            15'b11100011_0011_010: DATA = 1'b0;
            15'b11100011_0011_011: DATA = 1'b0;
            15'b11100011_0011_100: DATA = 1'b0;
            15'b11100011_0011_101: DATA = 1'b0;
            15'b11100011_0011_110: DATA = 1'b0;
            15'b11100011_0011_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 1 Row 4
            15'b11100011_0100_000: DATA = 1'b0;
            15'b11100011_0100_001: DATA = 1'b0;
            15'b11100011_0100_010: DATA = 1'b0;
            15'b11100011_0100_011: DATA = 1'b0;
            15'b11100011_0100_100: DATA = 1'b0;
            15'b11100011_0100_101: DATA = 1'b0;
            15'b11100011_0100_110: DATA = 1'b0;
            15'b11100011_0100_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 1 Row 5
            15'b11100011_0101_000: DATA = 1'b0;
            15'b11100011_0101_001: DATA = 1'b0;
            15'b11100011_0101_010: DATA = 1'b0;
            15'b11100011_0101_011: DATA = 1'b0;
            15'b11100011_0101_100: DATA = 1'b0;
            15'b11100011_0101_101: DATA = 1'b0;
            15'b11100011_0101_110: DATA = 1'b0;
            15'b11100011_0101_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 1 Row 6
            15'b11100011_0110_000: DATA = 1'b1;
            15'b11100011_0110_001: DATA = 1'b0;
            15'b11100011_0110_010: DATA = 1'b0;
            15'b11100011_0110_011: DATA = 1'b0;
            15'b11100011_0110_100: DATA = 1'b0;
            15'b11100011_0110_101: DATA = 1'b0;
            15'b11100011_0110_110: DATA = 1'b0;
            15'b11100011_0110_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 1 Row 7
            15'b11100011_0111_000: DATA = 1'b1;
            15'b11100011_0111_001: DATA = 1'b1;
            15'b11100011_0111_010: DATA = 1'b1;
            15'b11100011_0111_011: DATA = 1'b0;
            15'b11100011_0111_100: DATA = 1'b0;
            15'b11100011_0111_101: DATA = 1'b0;
            15'b11100011_0111_110: DATA = 1'b0;
            15'b11100011_0111_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 1 Row 8
            15'b11100011_1000_000: DATA = 1'b0;
            15'b11100011_1000_001: DATA = 1'b0;
            15'b11100011_1000_010: DATA = 1'b1;
            15'b11100011_1000_011: DATA = 1'b1;
            15'b11100011_1000_100: DATA = 1'b0;
            15'b11100011_1000_101: DATA = 1'b0;
            15'b11100011_1000_110: DATA = 1'b0;
            15'b11100011_1000_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 1 Row 9
            15'b11100011_1001_000: DATA = 1'b0;
            15'b11100011_1001_001: DATA = 1'b0;
            15'b11100011_1001_010: DATA = 1'b0;
            15'b11100011_1001_011: DATA = 1'b1;
            15'b11100011_1001_100: DATA = 1'b1;
            15'b11100011_1001_101: DATA = 1'b0;
            15'b11100011_1001_110: DATA = 1'b0;
            15'b11100011_1001_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 1 Row 10
            15'b11100011_1010_000: DATA = 1'b0;
            15'b11100011_1010_001: DATA = 1'b0;
            15'b11100011_1010_010: DATA = 1'b0;
            15'b11100011_1010_011: DATA = 1'b0;
            15'b11100011_1010_100: DATA = 1'b1;
            15'b11100011_1010_101: DATA = 1'b1;
            15'b11100011_1010_110: DATA = 1'b0;
            15'b11100011_1010_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 1 Row 11
            15'b11100011_1011_000: DATA = 1'b0;
            15'b11100011_1011_001: DATA = 1'b0;
            15'b11100011_1011_010: DATA = 1'b0;
            15'b11100011_1011_011: DATA = 1'b0;
            15'b11100011_1011_100: DATA = 1'b0;
            15'b11100011_1011_101: DATA = 1'b1;
            15'b11100011_1011_110: DATA = 1'b1;
            15'b11100011_1011_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 0 COL 1 Row 12
            15'b11100011_1100_000: DATA = 1'b0;
            15'b11100011_1100_001: DATA = 1'b0;
            15'b11100011_1100_010: DATA = 1'b0;
            15'b11100011_1100_011: DATA = 1'b0;
            15'b11100011_1100_100: DATA = 1'b0;
            15'b11100011_1100_101: DATA = 1'b0;
            15'b11100011_1100_110: DATA = 1'b0;
            15'b11100011_1100_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 0 COL 1 Row 13
            15'b11100011_1101_000: DATA = 1'b0;
            15'b11100011_1101_001: DATA = 1'b0;
            15'b11100011_1101_010: DATA = 1'b0;
            15'b11100011_1101_011: DATA = 1'b0;
            15'b11100011_1101_100: DATA = 1'b0;
            15'b11100011_1101_101: DATA = 1'b0;
            15'b11100011_1101_110: DATA = 1'b0;
            15'b11100011_1101_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 1 Row 14
            15'b11100011_1110_000: DATA = 1'b0;
            15'b11100011_1110_001: DATA = 1'b0;
            15'b11100011_1110_010: DATA = 1'b0;
            15'b11100011_1110_011: DATA = 1'b0;
            15'b11100011_1110_100: DATA = 1'b0;
            15'b11100011_1110_101: DATA = 1'b0;
            15'b11100011_1110_110: DATA = 1'b0;
            15'b11100011_1110_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 1 Row 15
            15'b11100011_1111_000: DATA = 1'b0;
            15'b11100011_1111_001: DATA = 1'b0;
            15'b11100011_1111_010: DATA = 1'b0;
            15'b11100011_1111_011: DATA = 1'b0;
            15'b11100011_1111_100: DATA = 1'b0;
            15'b11100011_1111_101: DATA = 1'b0;
            15'b11100011_1111_110: DATA = 1'b0;
            15'b11100011_1111_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 2 Row 0
            15'b11100100_0000_000: DATA = 1'b0;
            15'b11100100_0000_001: DATA = 1'b0;
            15'b11100100_0000_010: DATA = 1'b0;
            15'b11100100_0000_011: DATA = 1'b0;
            15'b11100100_0000_100: DATA = 1'b0;
            15'b11100100_0000_101: DATA = 1'b0;
            15'b11100100_0000_110: DATA = 1'b0;
            15'b11100100_0000_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 2 Row 1
            15'b11100100_0001_000: DATA = 1'b0;
            15'b11100100_0001_001: DATA = 1'b0;
            15'b11100100_0001_010: DATA = 1'b0;
            15'b11100100_0001_011: DATA = 1'b0;
            15'b11100100_0001_100: DATA = 1'b0;
            15'b11100100_0001_101: DATA = 1'b0;
            15'b11100100_0001_110: DATA = 1'b0;
            15'b11100100_0001_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 2 Row 2
            15'b11100100_0010_000: DATA = 1'b0;
            15'b11100100_0010_001: DATA = 1'b0;
            15'b11100100_0010_010: DATA = 1'b0;
            15'b11100100_0010_011: DATA = 1'b0;
            15'b11100100_0010_100: DATA = 1'b0;
            15'b11100100_0010_101: DATA = 1'b0;
            15'b11100100_0010_110: DATA = 1'b0;
            15'b11100100_0010_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 2 Row 3
            15'b11100100_0011_000: DATA = 1'b0;
            15'b11100100_0011_001: DATA = 1'b0;
            15'b11100100_0011_010: DATA = 1'b0;
            15'b11100100_0011_011: DATA = 1'b0;
            15'b11100100_0011_100: DATA = 1'b0;
            15'b11100100_0011_101: DATA = 1'b0;
            15'b11100100_0011_110: DATA = 1'b0;
            15'b11100100_0011_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 2 Row 4
            15'b11100100_0100_000: DATA = 1'b0;
            15'b11100100_0100_001: DATA = 1'b0;
            15'b11100100_0100_010: DATA = 1'b0;
            15'b11100100_0100_011: DATA = 1'b0;
            15'b11100100_0100_100: DATA = 1'b0;
            15'b11100100_0100_101: DATA = 1'b0;
            15'b11100100_0100_110: DATA = 1'b0;
            15'b11100100_0100_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 2 Row 5
            15'b11100100_0101_000: DATA = 1'b0;
            15'b11100100_0101_001: DATA = 1'b0;
            15'b11100100_0101_010: DATA = 1'b0;
            15'b11100100_0101_011: DATA = 1'b0;
            15'b11100100_0101_100: DATA = 1'b0;
            15'b11100100_0101_101: DATA = 1'b0;
            15'b11100100_0101_110: DATA = 1'b0;
            15'b11100100_0101_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 2 Row 6
            15'b11100100_0110_000: DATA = 1'b0;
            15'b11100100_0110_001: DATA = 1'b0;
            15'b11100100_0110_010: DATA = 1'b0;
            15'b11100100_0110_011: DATA = 1'b0;
            15'b11100100_0110_100: DATA = 1'b0;
            15'b11100100_0110_101: DATA = 1'b0;
            15'b11100100_0110_110: DATA = 1'b0;
            15'b11100100_0110_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 2 Row 7
            15'b11100100_0111_000: DATA = 1'b0;
            15'b11100100_0111_001: DATA = 1'b0;
            15'b11100100_0111_010: DATA = 1'b0;
            15'b11100100_0111_011: DATA = 1'b0;
            15'b11100100_0111_100: DATA = 1'b0;
            15'b11100100_0111_101: DATA = 1'b0;
            15'b11100100_0111_110: DATA = 1'b0;
            15'b11100100_0111_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 2 Row 8
            15'b11100100_1000_000: DATA = 1'b0;
            15'b11100100_1000_001: DATA = 1'b0;
            15'b11100100_1000_010: DATA = 1'b0;
            15'b11100100_1000_011: DATA = 1'b0;
            15'b11100100_1000_100: DATA = 1'b0;
            15'b11100100_1000_101: DATA = 1'b0;
            15'b11100100_1000_110: DATA = 1'b0;
            15'b11100100_1000_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 2 Row 9
            15'b11100100_1001_000: DATA = 1'b0;
            15'b11100100_1001_001: DATA = 1'b0;
            15'b11100100_1001_010: DATA = 1'b0;
            15'b11100100_1001_011: DATA = 1'b0;
            15'b11100100_1001_100: DATA = 1'b0;
            15'b11100100_1001_101: DATA = 1'b0;
            15'b11100100_1001_110: DATA = 1'b0;
            15'b11100100_1001_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 2 Row 10
            15'b11100100_1010_000: DATA = 1'b0;
            15'b11100100_1010_001: DATA = 1'b0;
            15'b11100100_1010_010: DATA = 1'b0;
            15'b11100100_1010_011: DATA = 1'b0;
            15'b11100100_1010_100: DATA = 1'b0;
            15'b11100100_1010_101: DATA = 1'b0;
            15'b11100100_1010_110: DATA = 1'b0;
            15'b11100100_1010_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 2 Row 11
            15'b11100100_1011_000: DATA = 1'b0;
            15'b11100100_1011_001: DATA = 1'b0;
            15'b11100100_1011_010: DATA = 1'b0;
            15'b11100100_1011_011: DATA = 1'b0;
            15'b11100100_1011_100: DATA = 1'b0;
            15'b11100100_1011_101: DATA = 1'b0;
            15'b11100100_1011_110: DATA = 1'b0;
            15'b11100100_1011_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 2 Row 12
            15'b11100100_1100_000: DATA = 1'b1;
            15'b11100100_1100_001: DATA = 1'b0;
            15'b11100100_1100_010: DATA = 1'b0;
            15'b11100100_1100_011: DATA = 1'b0;
            15'b11100100_1100_100: DATA = 1'b0;
            15'b11100100_1100_101: DATA = 1'b0;
            15'b11100100_1100_110: DATA = 1'b0;
            15'b11100100_1100_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 2 Row 13
            15'b11100100_1101_000: DATA = 1'b1;
            15'b11100100_1101_001: DATA = 1'b1;
            15'b11100100_1101_010: DATA = 1'b0;
            15'b11100100_1101_011: DATA = 1'b0;
            15'b11100100_1101_100: DATA = 1'b0;
            15'b11100100_1101_101: DATA = 1'b0;
            15'b11100100_1101_110: DATA = 1'b0;
            15'b11100100_1101_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 2 Row 14
            15'b11100100_1110_000: DATA = 1'b0;
            15'b11100100_1110_001: DATA = 1'b1;
            15'b11100100_1110_010: DATA = 1'b1;
            15'b11100100_1110_011: DATA = 1'b0;
            15'b11100100_1110_100: DATA = 1'b0;
            15'b11100100_1110_101: DATA = 1'b0;
            15'b11100100_1110_110: DATA = 1'b0;
            15'b11100100_1110_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 2 Row 15
            15'b11100100_1111_000: DATA = 1'b0;
            15'b11100100_1111_001: DATA = 1'b0;
            15'b11100100_1111_010: DATA = 1'b1;
            15'b11100100_1111_011: DATA = 1'b1;
            15'b11100100_1111_100: DATA = 1'b1;
            15'b11100100_1111_101: DATA = 1'b0;
            15'b11100100_1111_110: DATA = 1'b0;
            15'b11100100_1111_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 3 Row 0
            15'b11100101_0000_000: DATA = 1'b0;
            15'b11100101_0000_001: DATA = 1'b0;
            15'b11100101_0000_010: DATA = 1'b0;
            15'b11100101_0000_011: DATA = 1'b0;
            15'b11100101_0000_100: DATA = 1'b0;
            15'b11100101_0000_101: DATA = 1'b0;
            15'b11100101_0000_110: DATA = 1'b0;
            15'b11100101_0000_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 3 Row 1
            15'b11100101_0001_000: DATA = 1'b0;
            15'b11100101_0001_001: DATA = 1'b0;
            15'b11100101_0001_010: DATA = 1'b0;
            15'b11100101_0001_011: DATA = 1'b0;
            15'b11100101_0001_100: DATA = 1'b0;
            15'b11100101_0001_101: DATA = 1'b0;
            15'b11100101_0001_110: DATA = 1'b0;
            15'b11100101_0001_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 3 Row 2
            15'b11100101_0010_000: DATA = 1'b0;
            15'b11100101_0010_001: DATA = 1'b0;
            15'b11100101_0010_010: DATA = 1'b0;
            15'b11100101_0010_011: DATA = 1'b0;
            15'b11100101_0010_100: DATA = 1'b0;
            15'b11100101_0010_101: DATA = 1'b0;
            15'b11100101_0010_110: DATA = 1'b0;
            15'b11100101_0010_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 3 Row 3
            15'b11100101_0011_000: DATA = 1'b0;
            15'b11100101_0011_001: DATA = 1'b0;
            15'b11100101_0011_010: DATA = 1'b0;
            15'b11100101_0011_011: DATA = 1'b0;
            15'b11100101_0011_100: DATA = 1'b0;
            15'b11100101_0011_101: DATA = 1'b0;
            15'b11100101_0011_110: DATA = 1'b0;
            15'b11100101_0011_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 3 Row 4
            15'b11100101_0100_000: DATA = 1'b0;
            15'b11100101_0100_001: DATA = 1'b0;
            15'b11100101_0100_010: DATA = 1'b0;
            15'b11100101_0100_011: DATA = 1'b0;
            15'b11100101_0100_100: DATA = 1'b0;
            15'b11100101_0100_101: DATA = 1'b0;
            15'b11100101_0100_110: DATA = 1'b0;
            15'b11100101_0100_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 3 Row 5
            15'b11100101_0101_000: DATA = 1'b0;
            15'b11100101_0101_001: DATA = 1'b0;
            15'b11100101_0101_010: DATA = 1'b0;
            15'b11100101_0101_011: DATA = 1'b0;
            15'b11100101_0101_100: DATA = 1'b0;
            15'b11100101_0101_101: DATA = 1'b0;
            15'b11100101_0101_110: DATA = 1'b0;
            15'b11100101_0101_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 3 Row 6
            15'b11100101_0110_000: DATA = 1'b0;
            15'b11100101_0110_001: DATA = 1'b0;
            15'b11100101_0110_010: DATA = 1'b0;
            15'b11100101_0110_011: DATA = 1'b0;
            15'b11100101_0110_100: DATA = 1'b0;
            15'b11100101_0110_101: DATA = 1'b0;
            15'b11100101_0110_110: DATA = 1'b0;
            15'b11100101_0110_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 3 Row 7
            15'b11100101_0111_000: DATA = 1'b0;
            15'b11100101_0111_001: DATA = 1'b0;
            15'b11100101_0111_010: DATA = 1'b0;
            15'b11100101_0111_011: DATA = 1'b0;
            15'b11100101_0111_100: DATA = 1'b0;
            15'b11100101_0111_101: DATA = 1'b0;
            15'b11100101_0111_110: DATA = 1'b0;
            15'b11100101_0111_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 3 Row 8
            15'b11100101_1000_000: DATA = 1'b0;
            15'b11100101_1000_001: DATA = 1'b0;
            15'b11100101_1000_010: DATA = 1'b0;
            15'b11100101_1000_011: DATA = 1'b0;
            15'b11100101_1000_100: DATA = 1'b0;
            15'b11100101_1000_101: DATA = 1'b0;
            15'b11100101_1000_110: DATA = 1'b0;
            15'b11100101_1000_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 3 Row 9
            15'b11100101_1001_000: DATA = 1'b0;
            15'b11100101_1001_001: DATA = 1'b0;
            15'b11100101_1001_010: DATA = 1'b0;
            15'b11100101_1001_011: DATA = 1'b0;
            15'b11100101_1001_100: DATA = 1'b0;
            15'b11100101_1001_101: DATA = 1'b0;
            15'b11100101_1001_110: DATA = 1'b0;
            15'b11100101_1001_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 3 Row 10
            15'b11100101_1010_000: DATA = 1'b0;
            15'b11100101_1010_001: DATA = 1'b0;
            15'b11100101_1010_010: DATA = 1'b0;
            15'b11100101_1010_011: DATA = 1'b0;
            15'b11100101_1010_100: DATA = 1'b0;
            15'b11100101_1010_101: DATA = 1'b0;
            15'b11100101_1010_110: DATA = 1'b0;
            15'b11100101_1010_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 3 Row 11
            15'b11100101_1011_000: DATA = 1'b0;
            15'b11100101_1011_001: DATA = 1'b0;
            15'b11100101_1011_010: DATA = 1'b0;
            15'b11100101_1011_011: DATA = 1'b0;
            15'b11100101_1011_100: DATA = 1'b0;
            15'b11100101_1011_101: DATA = 1'b0;
            15'b11100101_1011_110: DATA = 1'b0;
            15'b11100101_1011_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 3 Row 12
            15'b11100101_1100_000: DATA = 1'b0;
            15'b11100101_1100_001: DATA = 1'b0;
            15'b11100101_1100_010: DATA = 1'b0;
            15'b11100101_1100_011: DATA = 1'b0;
            15'b11100101_1100_100: DATA = 1'b0;
            15'b11100101_1100_101: DATA = 1'b0;
            15'b11100101_1100_110: DATA = 1'b0;
            15'b11100101_1100_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 3 Row 13
            15'b11100101_1101_000: DATA = 1'b0;
            15'b11100101_1101_001: DATA = 1'b0;
            15'b11100101_1101_010: DATA = 1'b0;
            15'b11100101_1101_011: DATA = 1'b0;
            15'b11100101_1101_100: DATA = 1'b0;
            15'b11100101_1101_101: DATA = 1'b0;
            15'b11100101_1101_110: DATA = 1'b0;
            15'b11100101_1101_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 3 Row 14
            15'b11100101_1110_000: DATA = 1'b0;
            15'b11100101_1110_001: DATA = 1'b0;
            15'b11100101_1110_010: DATA = 1'b0;
            15'b11100101_1110_011: DATA = 1'b0;
            15'b11100101_1110_100: DATA = 1'b0;
            15'b11100101_1110_101: DATA = 1'b0;
            15'b11100101_1110_110: DATA = 1'b0;
            15'b11100101_1110_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 3 Row 15
            15'b11100101_1111_000: DATA = 1'b0;
            15'b11100101_1111_001: DATA = 1'b0;
            15'b11100101_1111_010: DATA = 1'b0;
            15'b11100101_1111_011: DATA = 1'b0;
            15'b11100101_1111_100: DATA = 1'b0;
            15'b11100101_1111_101: DATA = 1'b0;
            15'b11100101_1111_110: DATA = 1'b0;
            15'b11100101_1111_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 0 COL 4 Row 0
            15'b11100110_0000_000: DATA = 1'b0;
            15'b11100110_0000_001: DATA = 1'b0;
            15'b11100110_0000_010: DATA = 1'b0;
            15'b11100110_0000_011: DATA = 1'b0;
            15'b11100110_0000_100: DATA = 1'b0;
            15'b11100110_0000_101: DATA = 1'b0;
            15'b11100110_0000_110: DATA = 1'b0;
            15'b11100110_0000_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 0 COL 4 Row 1
            15'b11100110_0001_000: DATA = 1'b0;
            15'b11100110_0001_001: DATA = 1'b0;
            15'b11100110_0001_010: DATA = 1'b0;
            15'b11100110_0001_011: DATA = 1'b0;
            15'b11100110_0001_100: DATA = 1'b0;
            15'b11100110_0001_101: DATA = 1'b0;
            15'b11100110_0001_110: DATA = 1'b0;
            15'b11100110_0001_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 0 COL 4 Row 2
            15'b11100110_0010_000: DATA = 1'b0;
            15'b11100110_0010_001: DATA = 1'b0;
            15'b11100110_0010_010: DATA = 1'b0;
            15'b11100110_0010_011: DATA = 1'b0;
            15'b11100110_0010_100: DATA = 1'b0;
            15'b11100110_0010_101: DATA = 1'b0;
            15'b11100110_0010_110: DATA = 1'b0;
            15'b11100110_0010_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 0 COL 4 Row 3
            15'b11100110_0011_000: DATA = 1'b0;
            15'b11100110_0011_001: DATA = 1'b0;
            15'b11100110_0011_010: DATA = 1'b0;
            15'b11100110_0011_011: DATA = 1'b0;
            15'b11100110_0011_100: DATA = 1'b0;
            15'b11100110_0011_101: DATA = 1'b0;
            15'b11100110_0011_110: DATA = 1'b0;
            15'b11100110_0011_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 0 COL 4 Row 4
            15'b11100110_0100_000: DATA = 1'b0;
            15'b11100110_0100_001: DATA = 1'b0;
            15'b11100110_0100_010: DATA = 1'b0;
            15'b11100110_0100_011: DATA = 1'b0;
            15'b11100110_0100_100: DATA = 1'b0;
            15'b11100110_0100_101: DATA = 1'b0;
            15'b11100110_0100_110: DATA = 1'b0;
            15'b11100110_0100_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 0 COL 4 Row 5
            15'b11100110_0101_000: DATA = 1'b0;
            15'b11100110_0101_001: DATA = 1'b0;
            15'b11100110_0101_010: DATA = 1'b0;
            15'b11100110_0101_011: DATA = 1'b0;
            15'b11100110_0101_100: DATA = 1'b0;
            15'b11100110_0101_101: DATA = 1'b0;
            15'b11100110_0101_110: DATA = 1'b0;
            15'b11100110_0101_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 0 COL 4 Row 6
            15'b11100110_0110_000: DATA = 1'b0;
            15'b11100110_0110_001: DATA = 1'b0;
            15'b11100110_0110_010: DATA = 1'b0;
            15'b11100110_0110_011: DATA = 1'b0;
            15'b11100110_0110_100: DATA = 1'b0;
            15'b11100110_0110_101: DATA = 1'b0;
            15'b11100110_0110_110: DATA = 1'b0;
            15'b11100110_0110_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 0 COL 4 Row 7
            15'b11100110_0111_000: DATA = 1'b0;
            15'b11100110_0111_001: DATA = 1'b0;
            15'b11100110_0111_010: DATA = 1'b0;
            15'b11100110_0111_011: DATA = 1'b0;
            15'b11100110_0111_100: DATA = 1'b0;
            15'b11100110_0111_101: DATA = 1'b0;
            15'b11100110_0111_110: DATA = 1'b0;
            15'b11100110_0111_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 0 COL 4 Row 8
            15'b11100110_1000_000: DATA = 1'b0;
            15'b11100110_1000_001: DATA = 1'b0;
            15'b11100110_1000_010: DATA = 1'b0;
            15'b11100110_1000_011: DATA = 1'b0;
            15'b11100110_1000_100: DATA = 1'b0;
            15'b11100110_1000_101: DATA = 1'b0;
            15'b11100110_1000_110: DATA = 1'b0;
            15'b11100110_1000_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 0 COL 4 Row 9
            15'b11100110_1001_000: DATA = 1'b0;
            15'b11100110_1001_001: DATA = 1'b0;
            15'b11100110_1001_010: DATA = 1'b0;
            15'b11100110_1001_011: DATA = 1'b0;
            15'b11100110_1001_100: DATA = 1'b0;
            15'b11100110_1001_101: DATA = 1'b0;
            15'b11100110_1001_110: DATA = 1'b0;
            15'b11100110_1001_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 0 COL 4 Row 10
            15'b11100110_1010_000: DATA = 1'b0;
            15'b11100110_1010_001: DATA = 1'b0;
            15'b11100110_1010_010: DATA = 1'b0;
            15'b11100110_1010_011: DATA = 1'b0;
            15'b11100110_1010_100: DATA = 1'b0;
            15'b11100110_1010_101: DATA = 1'b0;
            15'b11100110_1010_110: DATA = 1'b0;
            15'b11100110_1010_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 0 COL 4 Row 11
            15'b11100110_1011_000: DATA = 1'b0;
            15'b11100110_1011_001: DATA = 1'b0;
            15'b11100110_1011_010: DATA = 1'b0;
            15'b11100110_1011_011: DATA = 1'b0;
            15'b11100110_1011_100: DATA = 1'b0;
            15'b11100110_1011_101: DATA = 1'b0;
            15'b11100110_1011_110: DATA = 1'b0;
            15'b11100110_1011_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 0 COL 4 Row 12
            15'b11100110_1100_000: DATA = 1'b0;
            15'b11100110_1100_001: DATA = 1'b0;
            15'b11100110_1100_010: DATA = 1'b0;
            15'b11100110_1100_011: DATA = 1'b0;
            15'b11100110_1100_100: DATA = 1'b0;
            15'b11100110_1100_101: DATA = 1'b0;
            15'b11100110_1100_110: DATA = 1'b0;
            15'b11100110_1100_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 0 COL 4 Row 13
            15'b11100110_1101_000: DATA = 1'b0;
            15'b11100110_1101_001: DATA = 1'b0;
            15'b11100110_1101_010: DATA = 1'b0;
            15'b11100110_1101_011: DATA = 1'b0;
            15'b11100110_1101_100: DATA = 1'b0;
            15'b11100110_1101_101: DATA = 1'b0;
            15'b11100110_1101_110: DATA = 1'b0;
            15'b11100110_1101_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 0 COL 4 Row 14
            15'b11100110_1110_000: DATA = 1'b0;
            15'b11100110_1110_001: DATA = 1'b0;
            15'b11100110_1110_010: DATA = 1'b0;
            15'b11100110_1110_011: DATA = 1'b0;
            15'b11100110_1110_100: DATA = 1'b0;
            15'b11100110_1110_101: DATA = 1'b0;
            15'b11100110_1110_110: DATA = 1'b0;
            15'b11100110_1110_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 0 COL 4 Row 15
            15'b11100110_1111_000: DATA = 1'b0;
            15'b11100110_1111_001: DATA = 1'b0;
            15'b11100110_1111_010: DATA = 1'b0;
            15'b11100110_1111_011: DATA = 1'b0;
            15'b11100110_1111_100: DATA = 1'b0;
            15'b11100110_1111_101: DATA = 1'b0;
            15'b11100110_1111_110: DATA = 1'b0;
            15'b11100110_1111_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 1 COL 0 Row 0
            15'b11100111_0000_000: DATA = 1'b0;
            15'b11100111_0000_001: DATA = 1'b0;
            15'b11100111_0000_010: DATA = 1'b0;
            15'b11100111_0000_011: DATA = 1'b0;
            15'b11100111_0000_100: DATA = 1'b0;
            15'b11100111_0000_101: DATA = 1'b0;
            15'b11100111_0000_110: DATA = 1'b0;
            15'b11100111_0000_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 0 Row 1
            15'b11100111_0001_000: DATA = 1'b0;
            15'b11100111_0001_001: DATA = 1'b0;
            15'b11100111_0001_010: DATA = 1'b0;
            15'b11100111_0001_011: DATA = 1'b0;
            15'b11100111_0001_100: DATA = 1'b0;
            15'b11100111_0001_101: DATA = 1'b0;
            15'b11100111_0001_110: DATA = 1'b0;
            15'b11100111_0001_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 0 Row 2
            15'b11100111_0010_000: DATA = 1'b0;
            15'b11100111_0010_001: DATA = 1'b0;
            15'b11100111_0010_010: DATA = 1'b0;
            15'b11100111_0010_011: DATA = 1'b0;
            15'b11100111_0010_100: DATA = 1'b0;
            15'b11100111_0010_101: DATA = 1'b0;
            15'b11100111_0010_110: DATA = 1'b0;
            15'b11100111_0010_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 0 Row 3
            15'b11100111_0011_000: DATA = 1'b0;
            15'b11100111_0011_001: DATA = 1'b0;
            15'b11100111_0011_010: DATA = 1'b0;
            15'b11100111_0011_011: DATA = 1'b0;
            15'b11100111_0011_100: DATA = 1'b0;
            15'b11100111_0011_101: DATA = 1'b0;
            15'b11100111_0011_110: DATA = 1'b0;
            15'b11100111_0011_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 0 Row 4
            15'b11100111_0100_000: DATA = 1'b0;
            15'b11100111_0100_001: DATA = 1'b0;
            15'b11100111_0100_010: DATA = 1'b0;
            15'b11100111_0100_011: DATA = 1'b0;
            15'b11100111_0100_100: DATA = 1'b0;
            15'b11100111_0100_101: DATA = 1'b0;
            15'b11100111_0100_110: DATA = 1'b0;
            15'b11100111_0100_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 0 Row 5
            15'b11100111_0101_000: DATA = 1'b0;
            15'b11100111_0101_001: DATA = 1'b0;
            15'b11100111_0101_010: DATA = 1'b0;
            15'b11100111_0101_011: DATA = 1'b0;
            15'b11100111_0101_100: DATA = 1'b0;
            15'b11100111_0101_101: DATA = 1'b0;
            15'b11100111_0101_110: DATA = 1'b0;
            15'b11100111_0101_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 0 Row 6
            15'b11100111_0110_000: DATA = 1'b0;
            15'b11100111_0110_001: DATA = 1'b0;
            15'b11100111_0110_010: DATA = 1'b0;
            15'b11100111_0110_011: DATA = 1'b0;
            15'b11100111_0110_100: DATA = 1'b0;
            15'b11100111_0110_101: DATA = 1'b0;
            15'b11100111_0110_110: DATA = 1'b0;
            15'b11100111_0110_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 0 Row 7
            15'b11100111_0111_000: DATA = 1'b0;
            15'b11100111_0111_001: DATA = 1'b0;
            15'b11100111_0111_010: DATA = 1'b0;
            15'b11100111_0111_011: DATA = 1'b0;
            15'b11100111_0111_100: DATA = 1'b0;
            15'b11100111_0111_101: DATA = 1'b0;
            15'b11100111_0111_110: DATA = 1'b0;
            15'b11100111_0111_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 0 Row 8
            15'b11100111_1000_000: DATA = 1'b0;
            15'b11100111_1000_001: DATA = 1'b0;
            15'b11100111_1000_010: DATA = 1'b0;
            15'b11100111_1000_011: DATA = 1'b0;
            15'b11100111_1000_100: DATA = 1'b0;
            15'b11100111_1000_101: DATA = 1'b0;
            15'b11100111_1000_110: DATA = 1'b0;
            15'b11100111_1000_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 0 Row 9
            15'b11100111_1001_000: DATA = 1'b0;
            15'b11100111_1001_001: DATA = 1'b0;
            15'b11100111_1001_010: DATA = 1'b0;
            15'b11100111_1001_011: DATA = 1'b0;
            15'b11100111_1001_100: DATA = 1'b0;
            15'b11100111_1001_101: DATA = 1'b0;
            15'b11100111_1001_110: DATA = 1'b0;
            15'b11100111_1001_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 0 Row 10
            15'b11100111_1010_000: DATA = 1'b0;
            15'b11100111_1010_001: DATA = 1'b0;
            15'b11100111_1010_010: DATA = 1'b0;
            15'b11100111_1010_011: DATA = 1'b0;
            15'b11100111_1010_100: DATA = 1'b0;
            15'b11100111_1010_101: DATA = 1'b0;
            15'b11100111_1010_110: DATA = 1'b0;
            15'b11100111_1010_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 0 Row 11
            15'b11100111_1011_000: DATA = 1'b0;
            15'b11100111_1011_001: DATA = 1'b0;
            15'b11100111_1011_010: DATA = 1'b0;
            15'b11100111_1011_011: DATA = 1'b0;
            15'b11100111_1011_100: DATA = 1'b0;
            15'b11100111_1011_101: DATA = 1'b0;
            15'b11100111_1011_110: DATA = 1'b0;
            15'b11100111_1011_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 0 Row 12
            15'b11100111_1100_000: DATA = 1'b0;
            15'b11100111_1100_001: DATA = 1'b0;
            15'b11100111_1100_010: DATA = 1'b0;
            15'b11100111_1100_011: DATA = 1'b0;
            15'b11100111_1100_100: DATA = 1'b0;
            15'b11100111_1100_101: DATA = 1'b0;
            15'b11100111_1100_110: DATA = 1'b0;
            15'b11100111_1100_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 0 Row 13
            15'b11100111_1101_000: DATA = 1'b0;
            15'b11100111_1101_001: DATA = 1'b0;
            15'b11100111_1101_010: DATA = 1'b0;
            15'b11100111_1101_011: DATA = 1'b0;
            15'b11100111_1101_100: DATA = 1'b0;
            15'b11100111_1101_101: DATA = 1'b0;
            15'b11100111_1101_110: DATA = 1'b0;
            15'b11100111_1101_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 0 Row 14
            15'b11100111_1110_000: DATA = 1'b0;
            15'b11100111_1110_001: DATA = 1'b0;
            15'b11100111_1110_010: DATA = 1'b0;
            15'b11100111_1110_011: DATA = 1'b0;
            15'b11100111_1110_100: DATA = 1'b0;
            15'b11100111_1110_101: DATA = 1'b0;
            15'b11100111_1110_110: DATA = 1'b0;
            15'b11100111_1110_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 0 Row 15
            15'b11100111_1111_000: DATA = 1'b0;
            15'b11100111_1111_001: DATA = 1'b0;
            15'b11100111_1111_010: DATA = 1'b0;
            15'b11100111_1111_011: DATA = 1'b0;
            15'b11100111_1111_100: DATA = 1'b0;
            15'b11100111_1111_101: DATA = 1'b0;
            15'b11100111_1111_110: DATA = 1'b0;
            15'b11100111_1111_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 1 Row 0
            15'b11101000_0000_000: DATA = 1'b0;
            15'b11101000_0000_001: DATA = 1'b0;
            15'b11101000_0000_010: DATA = 1'b0;
            15'b11101000_0000_011: DATA = 1'b0;
            15'b11101000_0000_100: DATA = 1'b0;
            15'b11101000_0000_101: DATA = 1'b0;
            15'b11101000_0000_110: DATA = 1'b0;
            15'b11101000_0000_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 1 Row 1
            15'b11101000_0001_000: DATA = 1'b0;
            15'b11101000_0001_001: DATA = 1'b0;
            15'b11101000_0001_010: DATA = 1'b0;
            15'b11101000_0001_011: DATA = 1'b0;
            15'b11101000_0001_100: DATA = 1'b0;
            15'b11101000_0001_101: DATA = 1'b0;
            15'b11101000_0001_110: DATA = 1'b0;
            15'b11101000_0001_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 1 Row 2
            15'b11101000_0010_000: DATA = 1'b0;
            15'b11101000_0010_001: DATA = 1'b0;
            15'b11101000_0010_010: DATA = 1'b0;
            15'b11101000_0010_011: DATA = 1'b0;
            15'b11101000_0010_100: DATA = 1'b0;
            15'b11101000_0010_101: DATA = 1'b0;
            15'b11101000_0010_110: DATA = 1'b0;
            15'b11101000_0010_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 1 Row 3
            15'b11101000_0011_000: DATA = 1'b0;
            15'b11101000_0011_001: DATA = 1'b0;
            15'b11101000_0011_010: DATA = 1'b0;
            15'b11101000_0011_011: DATA = 1'b0;
            15'b11101000_0011_100: DATA = 1'b0;
            15'b11101000_0011_101: DATA = 1'b0;
            15'b11101000_0011_110: DATA = 1'b0;
            15'b11101000_0011_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 1 Row 4
            15'b11101000_0100_000: DATA = 1'b0;
            15'b11101000_0100_001: DATA = 1'b0;
            15'b11101000_0100_010: DATA = 1'b0;
            15'b11101000_0100_011: DATA = 1'b0;
            15'b11101000_0100_100: DATA = 1'b0;
            15'b11101000_0100_101: DATA = 1'b0;
            15'b11101000_0100_110: DATA = 1'b0;
            15'b11101000_0100_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 1 Row 5
            15'b11101000_0101_000: DATA = 1'b0;
            15'b11101000_0101_001: DATA = 1'b0;
            15'b11101000_0101_010: DATA = 1'b0;
            15'b11101000_0101_011: DATA = 1'b0;
            15'b11101000_0101_100: DATA = 1'b0;
            15'b11101000_0101_101: DATA = 1'b0;
            15'b11101000_0101_110: DATA = 1'b0;
            15'b11101000_0101_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 1 Row 6
            15'b11101000_0110_000: DATA = 1'b0;
            15'b11101000_0110_001: DATA = 1'b0;
            15'b11101000_0110_010: DATA = 1'b0;
            15'b11101000_0110_011: DATA = 1'b0;
            15'b11101000_0110_100: DATA = 1'b0;
            15'b11101000_0110_101: DATA = 1'b0;
            15'b11101000_0110_110: DATA = 1'b0;
            15'b11101000_0110_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 1 Row 7
            15'b11101000_0111_000: DATA = 1'b0;
            15'b11101000_0111_001: DATA = 1'b0;
            15'b11101000_0111_010: DATA = 1'b0;
            15'b11101000_0111_011: DATA = 1'b0;
            15'b11101000_0111_100: DATA = 1'b0;
            15'b11101000_0111_101: DATA = 1'b0;
            15'b11101000_0111_110: DATA = 1'b0;
            15'b11101000_0111_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 1 Row 8
            15'b11101000_1000_000: DATA = 1'b0;
            15'b11101000_1000_001: DATA = 1'b0;
            15'b11101000_1000_010: DATA = 1'b0;
            15'b11101000_1000_011: DATA = 1'b0;
            15'b11101000_1000_100: DATA = 1'b0;
            15'b11101000_1000_101: DATA = 1'b0;
            15'b11101000_1000_110: DATA = 1'b0;
            15'b11101000_1000_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 1 Row 9
            15'b11101000_1001_000: DATA = 1'b0;
            15'b11101000_1001_001: DATA = 1'b0;
            15'b11101000_1001_010: DATA = 1'b0;
            15'b11101000_1001_011: DATA = 1'b0;
            15'b11101000_1001_100: DATA = 1'b0;
            15'b11101000_1001_101: DATA = 1'b0;
            15'b11101000_1001_110: DATA = 1'b0;
            15'b11101000_1001_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 1 Row 10
            15'b11101000_1010_000: DATA = 1'b0;
            15'b11101000_1010_001: DATA = 1'b0;
            15'b11101000_1010_010: DATA = 1'b0;
            15'b11101000_1010_011: DATA = 1'b0;
            15'b11101000_1010_100: DATA = 1'b0;
            15'b11101000_1010_101: DATA = 1'b0;
            15'b11101000_1010_110: DATA = 1'b0;
            15'b11101000_1010_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 1 Row 11
            15'b11101000_1011_000: DATA = 1'b0;
            15'b11101000_1011_001: DATA = 1'b0;
            15'b11101000_1011_010: DATA = 1'b0;
            15'b11101000_1011_011: DATA = 1'b0;
            15'b11101000_1011_100: DATA = 1'b0;
            15'b11101000_1011_101: DATA = 1'b0;
            15'b11101000_1011_110: DATA = 1'b0;
            15'b11101000_1011_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 1 Row 12
            15'b11101000_1100_000: DATA = 1'b0;
            15'b11101000_1100_001: DATA = 1'b0;
            15'b11101000_1100_010: DATA = 1'b0;
            15'b11101000_1100_011: DATA = 1'b0;
            15'b11101000_1100_100: DATA = 1'b0;
            15'b11101000_1100_101: DATA = 1'b0;
            15'b11101000_1100_110: DATA = 1'b0;
            15'b11101000_1100_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 1 Row 13
            15'b11101000_1101_000: DATA = 1'b0;
            15'b11101000_1101_001: DATA = 1'b0;
            15'b11101000_1101_010: DATA = 1'b0;
            15'b11101000_1101_011: DATA = 1'b0;
            15'b11101000_1101_100: DATA = 1'b0;
            15'b11101000_1101_101: DATA = 1'b0;
            15'b11101000_1101_110: DATA = 1'b0;
            15'b11101000_1101_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 1 Row 14
            15'b11101000_1110_000: DATA = 1'b0;
            15'b11101000_1110_001: DATA = 1'b0;
            15'b11101000_1110_010: DATA = 1'b0;
            15'b11101000_1110_011: DATA = 1'b0;
            15'b11101000_1110_100: DATA = 1'b0;
            15'b11101000_1110_101: DATA = 1'b0;
            15'b11101000_1110_110: DATA = 1'b0;
            15'b11101000_1110_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 1 Row 15
            15'b11101000_1111_000: DATA = 1'b0;
            15'b11101000_1111_001: DATA = 1'b0;
            15'b11101000_1111_010: DATA = 1'b0;
            15'b11101000_1111_011: DATA = 1'b0;
            15'b11101000_1111_100: DATA = 1'b0;
            15'b11101000_1111_101: DATA = 1'b0;
            15'b11101000_1111_110: DATA = 1'b0;
            15'b11101000_1111_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 2 Row 0
            15'b11101001_0000_000: DATA = 1'b0;
            15'b11101001_0000_001: DATA = 1'b0;
            15'b11101001_0000_010: DATA = 1'b0;
            15'b11101001_0000_011: DATA = 1'b0;
            15'b11101001_0000_100: DATA = 1'b1;
            15'b11101001_0000_101: DATA = 1'b1;
            15'b11101001_0000_110: DATA = 1'b0;
            15'b11101001_0000_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 2 Row 1
            15'b11101001_0001_000: DATA = 1'b0;
            15'b11101001_0001_001: DATA = 1'b0;
            15'b11101001_0001_010: DATA = 1'b0;
            15'b11101001_0001_011: DATA = 1'b0;
            15'b11101001_0001_100: DATA = 1'b0;
            15'b11101001_0001_101: DATA = 1'b1;
            15'b11101001_0001_110: DATA = 1'b1;
            15'b11101001_0001_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 2 Row 2
            15'b11101001_0010_000: DATA = 1'b0;
            15'b11101001_0010_001: DATA = 1'b0;
            15'b11101001_0010_010: DATA = 1'b0;
            15'b11101001_0010_011: DATA = 1'b0;
            15'b11101001_0010_100: DATA = 1'b0;
            15'b11101001_0010_101: DATA = 1'b0;
            15'b11101001_0010_110: DATA = 1'b1;
            15'b11101001_0010_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 1 COL 2 Row 3
            15'b11101001_0011_000: DATA = 1'b0;
            15'b11101001_0011_001: DATA = 1'b0;
            15'b11101001_0011_010: DATA = 1'b0;
            15'b11101001_0011_011: DATA = 1'b0;
            15'b11101001_0011_100: DATA = 1'b0;
            15'b11101001_0011_101: DATA = 1'b0;
            15'b11101001_0011_110: DATA = 1'b0;
            15'b11101001_0011_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 1 COL 2 Row 4
            15'b11101001_0100_000: DATA = 1'b0;
            15'b11101001_0100_001: DATA = 1'b0;
            15'b11101001_0100_010: DATA = 1'b0;
            15'b11101001_0100_011: DATA = 1'b0;
            15'b11101001_0100_100: DATA = 1'b0;
            15'b11101001_0100_101: DATA = 1'b0;
            15'b11101001_0100_110: DATA = 1'b0;
            15'b11101001_0100_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 2 Row 5
            15'b11101001_0101_000: DATA = 1'b0;
            15'b11101001_0101_001: DATA = 1'b0;
            15'b11101001_0101_010: DATA = 1'b0;
            15'b11101001_0101_011: DATA = 1'b0;
            15'b11101001_0101_100: DATA = 1'b0;
            15'b11101001_0101_101: DATA = 1'b0;
            15'b11101001_0101_110: DATA = 1'b0;
            15'b11101001_0101_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 2 Row 6
            15'b11101001_0110_000: DATA = 1'b0;
            15'b11101001_0110_001: DATA = 1'b0;
            15'b11101001_0110_010: DATA = 1'b0;
            15'b11101001_0110_011: DATA = 1'b0;
            15'b11101001_0110_100: DATA = 1'b0;
            15'b11101001_0110_101: DATA = 1'b0;
            15'b11101001_0110_110: DATA = 1'b0;
            15'b11101001_0110_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 2 Row 7
            15'b11101001_0111_000: DATA = 1'b0;
            15'b11101001_0111_001: DATA = 1'b0;
            15'b11101001_0111_010: DATA = 1'b0;
            15'b11101001_0111_011: DATA = 1'b0;
            15'b11101001_0111_100: DATA = 1'b0;
            15'b11101001_0111_101: DATA = 1'b0;
            15'b11101001_0111_110: DATA = 1'b0;
            15'b11101001_0111_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 2 Row 8
            15'b11101001_1000_000: DATA = 1'b0;
            15'b11101001_1000_001: DATA = 1'b0;
            15'b11101001_1000_010: DATA = 1'b0;
            15'b11101001_1000_011: DATA = 1'b0;
            15'b11101001_1000_100: DATA = 1'b0;
            15'b11101001_1000_101: DATA = 1'b0;
            15'b11101001_1000_110: DATA = 1'b0;
            15'b11101001_1000_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 2 Row 9
            15'b11101001_1001_000: DATA = 1'b0;
            15'b11101001_1001_001: DATA = 1'b0;
            15'b11101001_1001_010: DATA = 1'b0;
            15'b11101001_1001_011: DATA = 1'b0;
            15'b11101001_1001_100: DATA = 1'b0;
            15'b11101001_1001_101: DATA = 1'b0;
            15'b11101001_1001_110: DATA = 1'b0;
            15'b11101001_1001_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 2 Row 10
            15'b11101001_1010_000: DATA = 1'b0;
            15'b11101001_1010_001: DATA = 1'b0;
            15'b11101001_1010_010: DATA = 1'b0;
            15'b11101001_1010_011: DATA = 1'b0;
            15'b11101001_1010_100: DATA = 1'b0;
            15'b11101001_1010_101: DATA = 1'b0;
            15'b11101001_1010_110: DATA = 1'b0;
            15'b11101001_1010_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 2 Row 11
            15'b11101001_1011_000: DATA = 1'b0;
            15'b11101001_1011_001: DATA = 1'b0;
            15'b11101001_1011_010: DATA = 1'b0;
            15'b11101001_1011_011: DATA = 1'b0;
            15'b11101001_1011_100: DATA = 1'b0;
            15'b11101001_1011_101: DATA = 1'b0;
            15'b11101001_1011_110: DATA = 1'b0;
            15'b11101001_1011_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 2 Row 12
            15'b11101001_1100_000: DATA = 1'b0;
            15'b11101001_1100_001: DATA = 1'b0;
            15'b11101001_1100_010: DATA = 1'b0;
            15'b11101001_1100_011: DATA = 1'b0;
            15'b11101001_1100_100: DATA = 1'b0;
            15'b11101001_1100_101: DATA = 1'b0;
            15'b11101001_1100_110: DATA = 1'b0;
            15'b11101001_1100_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 2 Row 13
            15'b11101001_1101_000: DATA = 1'b0;
            15'b11101001_1101_001: DATA = 1'b0;
            15'b11101001_1101_010: DATA = 1'b0;
            15'b11101001_1101_011: DATA = 1'b0;
            15'b11101001_1101_100: DATA = 1'b0;
            15'b11101001_1101_101: DATA = 1'b0;
            15'b11101001_1101_110: DATA = 1'b0;
            15'b11101001_1101_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 2 Row 14
            15'b11101001_1110_000: DATA = 1'b0;
            15'b11101001_1110_001: DATA = 1'b0;
            15'b11101001_1110_010: DATA = 1'b0;
            15'b11101001_1110_011: DATA = 1'b0;
            15'b11101001_1110_100: DATA = 1'b0;
            15'b11101001_1110_101: DATA = 1'b0;
            15'b11101001_1110_110: DATA = 1'b0;
            15'b11101001_1110_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 2 Row 15
            15'b11101001_1111_000: DATA = 1'b0;
            15'b11101001_1111_001: DATA = 1'b0;
            15'b11101001_1111_010: DATA = 1'b0;
            15'b11101001_1111_011: DATA = 1'b0;
            15'b11101001_1111_100: DATA = 1'b0;
            15'b11101001_1111_101: DATA = 1'b0;
            15'b11101001_1111_110: DATA = 1'b0;
            15'b11101001_1111_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 3 Row 0
            15'b11101010_0000_000: DATA = 1'b0;
            15'b11101010_0000_001: DATA = 1'b0;
            15'b11101010_0000_010: DATA = 1'b0;
            15'b11101010_0000_011: DATA = 1'b0;
            15'b11101010_0000_100: DATA = 1'b0;
            15'b11101010_0000_101: DATA = 1'b0;
            15'b11101010_0000_110: DATA = 1'b0;
            15'b11101010_0000_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 3 Row 1
            15'b11101010_0001_000: DATA = 1'b0;
            15'b11101010_0001_001: DATA = 1'b0;
            15'b11101010_0001_010: DATA = 1'b0;
            15'b11101010_0001_011: DATA = 1'b0;
            15'b11101010_0001_100: DATA = 1'b0;
            15'b11101010_0001_101: DATA = 1'b0;
            15'b11101010_0001_110: DATA = 1'b0;
            15'b11101010_0001_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 3 Row 2
            15'b11101010_0010_000: DATA = 1'b0;
            15'b11101010_0010_001: DATA = 1'b0;
            15'b11101010_0010_010: DATA = 1'b0;
            15'b11101010_0010_011: DATA = 1'b0;
            15'b11101010_0010_100: DATA = 1'b0;
            15'b11101010_0010_101: DATA = 1'b0;
            15'b11101010_0010_110: DATA = 1'b0;
            15'b11101010_0010_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 3 Row 3
            15'b11101010_0011_000: DATA = 1'b1;
            15'b11101010_0011_001: DATA = 1'b1;
            15'b11101010_0011_010: DATA = 1'b0;
            15'b11101010_0011_011: DATA = 1'b0;
            15'b11101010_0011_100: DATA = 1'b0;
            15'b11101010_0011_101: DATA = 1'b0;
            15'b11101010_0011_110: DATA = 1'b0;
            15'b11101010_0011_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 3 Row 4
            15'b11101010_0100_000: DATA = 1'b0;
            15'b11101010_0100_001: DATA = 1'b1;
            15'b11101010_0100_010: DATA = 1'b1;
            15'b11101010_0100_011: DATA = 1'b0;
            15'b11101010_0100_100: DATA = 1'b0;
            15'b11101010_0100_101: DATA = 1'b0;
            15'b11101010_0100_110: DATA = 1'b0;
            15'b11101010_0100_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 3 Row 5
            15'b11101010_0101_000: DATA = 1'b0;
            15'b11101010_0101_001: DATA = 1'b0;
            15'b11101010_0101_010: DATA = 1'b1;
            15'b11101010_0101_011: DATA = 1'b1;
            15'b11101010_0101_100: DATA = 1'b0;
            15'b11101010_0101_101: DATA = 1'b0;
            15'b11101010_0101_110: DATA = 1'b0;
            15'b11101010_0101_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 3 Row 6
            15'b11101010_0110_000: DATA = 1'b0;
            15'b11101010_0110_001: DATA = 1'b0;
            15'b11101010_0110_010: DATA = 1'b0;
            15'b11101010_0110_011: DATA = 1'b1;
            15'b11101010_0110_100: DATA = 1'b1;
            15'b11101010_0110_101: DATA = 1'b0;
            15'b11101010_0110_110: DATA = 1'b0;
            15'b11101010_0110_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 3 Row 7
            15'b11101010_0111_000: DATA = 1'b0;
            15'b11101010_0111_001: DATA = 1'b0;
            15'b11101010_0111_010: DATA = 1'b0;
            15'b11101010_0111_011: DATA = 1'b0;
            15'b11101010_0111_100: DATA = 1'b1;
            15'b11101010_0111_101: DATA = 1'b1;
            15'b11101010_0111_110: DATA = 1'b1;
            15'b11101010_0111_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 3 Row 8
            15'b11101010_1000_000: DATA = 1'b0;
            15'b11101010_1000_001: DATA = 1'b0;
            15'b11101010_1000_010: DATA = 1'b0;
            15'b11101010_1000_011: DATA = 1'b0;
            15'b11101010_1000_100: DATA = 1'b0;
            15'b11101010_1000_101: DATA = 1'b0;
            15'b11101010_1000_110: DATA = 1'b1;
            15'b11101010_1000_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 1 COL 3 Row 9
            15'b11101010_1001_000: DATA = 1'b0;
            15'b11101010_1001_001: DATA = 1'b0;
            15'b11101010_1001_010: DATA = 1'b0;
            15'b11101010_1001_011: DATA = 1'b0;
            15'b11101010_1001_100: DATA = 1'b0;
            15'b11101010_1001_101: DATA = 1'b0;
            15'b11101010_1001_110: DATA = 1'b0;
            15'b11101010_1001_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 1 COL 3 Row 10
            15'b11101010_1010_000: DATA = 1'b0;
            15'b11101010_1010_001: DATA = 1'b0;
            15'b11101010_1010_010: DATA = 1'b0;
            15'b11101010_1010_011: DATA = 1'b0;
            15'b11101010_1010_100: DATA = 1'b0;
            15'b11101010_1010_101: DATA = 1'b0;
            15'b11101010_1010_110: DATA = 1'b0;
            15'b11101010_1010_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 3 Row 11
            15'b11101010_1011_000: DATA = 1'b0;
            15'b11101010_1011_001: DATA = 1'b0;
            15'b11101010_1011_010: DATA = 1'b0;
            15'b11101010_1011_011: DATA = 1'b0;
            15'b11101010_1011_100: DATA = 1'b0;
            15'b11101010_1011_101: DATA = 1'b0;
            15'b11101010_1011_110: DATA = 1'b0;
            15'b11101010_1011_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 3 Row 12
            15'b11101010_1100_000: DATA = 1'b0;
            15'b11101010_1100_001: DATA = 1'b0;
            15'b11101010_1100_010: DATA = 1'b0;
            15'b11101010_1100_011: DATA = 1'b0;
            15'b11101010_1100_100: DATA = 1'b0;
            15'b11101010_1100_101: DATA = 1'b0;
            15'b11101010_1100_110: DATA = 1'b0;
            15'b11101010_1100_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 3 Row 13
            15'b11101010_1101_000: DATA = 1'b0;
            15'b11101010_1101_001: DATA = 1'b0;
            15'b11101010_1101_010: DATA = 1'b0;
            15'b11101010_1101_011: DATA = 1'b0;
            15'b11101010_1101_100: DATA = 1'b0;
            15'b11101010_1101_101: DATA = 1'b0;
            15'b11101010_1101_110: DATA = 1'b0;
            15'b11101010_1101_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 3 Row 14
            15'b11101010_1110_000: DATA = 1'b0;
            15'b11101010_1110_001: DATA = 1'b0;
            15'b11101010_1110_010: DATA = 1'b0;
            15'b11101010_1110_011: DATA = 1'b0;
            15'b11101010_1110_100: DATA = 1'b0;
            15'b11101010_1110_101: DATA = 1'b0;
            15'b11101010_1110_110: DATA = 1'b0;
            15'b11101010_1110_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 3 Row 15
            15'b11101010_1111_000: DATA = 1'b0;
            15'b11101010_1111_001: DATA = 1'b0;
            15'b11101010_1111_010: DATA = 1'b0;
            15'b11101010_1111_011: DATA = 1'b0;
            15'b11101010_1111_100: DATA = 1'b0;
            15'b11101010_1111_101: DATA = 1'b0;
            15'b11101010_1111_110: DATA = 1'b0;
            15'b11101010_1111_111: DATA = 1'b0;
            //SAWTOOTHY- ROW 1 COL 4 Row 0
            15'b11101011_0000_000: DATA = 1'b0;
            15'b11101011_0000_001: DATA = 1'b0;
            15'b11101011_0000_010: DATA = 1'b0;
            15'b11101011_0000_011: DATA = 1'b0;
            15'b11101011_0000_100: DATA = 1'b0;
            15'b11101011_0000_101: DATA = 1'b0;
            15'b11101011_0000_110: DATA = 1'b0;
            15'b11101011_0000_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 1 COL 4 Row 1
            15'b11101011_0001_000: DATA = 1'b0;
            15'b11101011_0001_001: DATA = 1'b0;
            15'b11101011_0001_010: DATA = 1'b0;
            15'b11101011_0001_011: DATA = 1'b0;
            15'b11101011_0001_100: DATA = 1'b0;
            15'b11101011_0001_101: DATA = 1'b0;
            15'b11101011_0001_110: DATA = 1'b0;
            15'b11101011_0001_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 1 COL 4 Row 2
            15'b11101011_0010_000: DATA = 1'b0;
            15'b11101011_0010_001: DATA = 1'b0;
            15'b11101011_0010_010: DATA = 1'b0;
            15'b11101011_0010_011: DATA = 1'b0;
            15'b11101011_0010_100: DATA = 1'b0;
            15'b11101011_0010_101: DATA = 1'b0;
            15'b11101011_0010_110: DATA = 1'b0;
            15'b11101011_0010_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 1 COL 4 Row 3
            15'b11101011_0011_000: DATA = 1'b0;
            15'b11101011_0011_001: DATA = 1'b0;
            15'b11101011_0011_010: DATA = 1'b0;
            15'b11101011_0011_011: DATA = 1'b0;
            15'b11101011_0011_100: DATA = 1'b0;
            15'b11101011_0011_101: DATA = 1'b0;
            15'b11101011_0011_110: DATA = 1'b0;
            15'b11101011_0011_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 1 COL 4 Row 4
            15'b11101011_0100_000: DATA = 1'b0;
            15'b11101011_0100_001: DATA = 1'b0;
            15'b11101011_0100_010: DATA = 1'b0;
            15'b11101011_0100_011: DATA = 1'b0;
            15'b11101011_0100_100: DATA = 1'b0;
            15'b11101011_0100_101: DATA = 1'b0;
            15'b11101011_0100_110: DATA = 1'b0;
            15'b11101011_0100_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 1 COL 4 Row 5
            15'b11101011_0101_000: DATA = 1'b0;
            15'b11101011_0101_001: DATA = 1'b0;
            15'b11101011_0101_010: DATA = 1'b0;
            15'b11101011_0101_011: DATA = 1'b0;
            15'b11101011_0101_100: DATA = 1'b0;
            15'b11101011_0101_101: DATA = 1'b0;
            15'b11101011_0101_110: DATA = 1'b0;
            15'b11101011_0101_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 1 COL 4 Row 6
            15'b11101011_0110_000: DATA = 1'b0;
            15'b11101011_0110_001: DATA = 1'b0;
            15'b11101011_0110_010: DATA = 1'b0;
            15'b11101011_0110_011: DATA = 1'b0;
            15'b11101011_0110_100: DATA = 1'b0;
            15'b11101011_0110_101: DATA = 1'b0;
            15'b11101011_0110_110: DATA = 1'b0;
            15'b11101011_0110_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 1 COL 4 Row 7
            15'b11101011_0111_000: DATA = 1'b0;
            15'b11101011_0111_001: DATA = 1'b0;
            15'b11101011_0111_010: DATA = 1'b0;
            15'b11101011_0111_011: DATA = 1'b0;
            15'b11101011_0111_100: DATA = 1'b0;
            15'b11101011_0111_101: DATA = 1'b0;
            15'b11101011_0111_110: DATA = 1'b0;
            15'b11101011_0111_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 1 COL 4 Row 8
            15'b11101011_1000_000: DATA = 1'b0;
            15'b11101011_1000_001: DATA = 1'b0;
            15'b11101011_1000_010: DATA = 1'b0;
            15'b11101011_1000_011: DATA = 1'b0;
            15'b11101011_1000_100: DATA = 1'b0;
            15'b11101011_1000_101: DATA = 1'b0;
            15'b11101011_1000_110: DATA = 1'b0;
            15'b11101011_1000_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 1 COL 4 Row 9
            15'b11101011_1001_000: DATA = 1'b1;
            15'b11101011_1001_001: DATA = 1'b0;
            15'b11101011_1001_010: DATA = 1'b0;
            15'b11101011_1001_011: DATA = 1'b0;
            15'b11101011_1001_100: DATA = 1'b0;
            15'b11101011_1001_101: DATA = 1'b0;
            15'b11101011_1001_110: DATA = 1'b0;
            15'b11101011_1001_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 1 COL 4 Row 10
            15'b11101011_1010_000: DATA = 1'b1;
            15'b11101011_1010_001: DATA = 1'b1;
            15'b11101011_1010_010: DATA = 1'b0;
            15'b11101011_1010_011: DATA = 1'b0;
            15'b11101011_1010_100: DATA = 1'b0;
            15'b11101011_1010_101: DATA = 1'b0;
            15'b11101011_1010_110: DATA = 1'b0;
            15'b11101011_1010_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 1 COL 4 Row 11
            15'b11101011_1011_000: DATA = 1'b0;
            15'b11101011_1011_001: DATA = 1'b1;
            15'b11101011_1011_010: DATA = 1'b1;
            15'b11101011_1011_011: DATA = 1'b1;
            15'b11101011_1011_100: DATA = 1'b0;
            15'b11101011_1011_101: DATA = 1'b0;
            15'b11101011_1011_110: DATA = 1'b0;
            15'b11101011_1011_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 1 COL 4 Row 12
            15'b11101011_1100_000: DATA = 1'b0;
            15'b11101011_1100_001: DATA = 1'b0;
            15'b11101011_1100_010: DATA = 1'b0;
            15'b11101011_1100_011: DATA = 1'b1;
            15'b11101011_1100_100: DATA = 1'b1;
            15'b11101011_1100_101: DATA = 1'b0;
            15'b11101011_1100_110: DATA = 1'b0;
            15'b11101011_1100_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 1 COL 4 Row 13
            15'b11101011_1101_000: DATA = 1'b0;
            15'b11101011_1101_001: DATA = 1'b0;
            15'b11101011_1101_010: DATA = 1'b0;
            15'b11101011_1101_011: DATA = 1'b0;
            15'b11101011_1101_100: DATA = 1'b1;
            15'b11101011_1101_101: DATA = 1'b1;
            15'b11101011_1101_110: DATA = 1'b0;
            15'b11101011_1101_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 1 COL 4 Row 14
            15'b11101011_1110_000: DATA = 1'b0;
            15'b11101011_1110_001: DATA = 1'b0;
            15'b11101011_1110_010: DATA = 1'b0;
            15'b11101011_1110_011: DATA = 1'b0;
            15'b11101011_1110_100: DATA = 1'b0;
            15'b11101011_1110_101: DATA = 1'b1;
            15'b11101011_1110_110: DATA = 1'b0;
            15'b11101011_1110_111: DATA = 1'b1;
            //SAWTOOTHY- ROW 1 COL 4 Row 15
            15'b11101011_1111_000: DATA = 1'b0;
            15'b11101011_1111_001: DATA = 1'b0;
            15'b11101011_1111_010: DATA = 1'b0;
            15'b11101011_1111_011: DATA = 1'b0;
            15'b11101011_1111_100: DATA = 1'b0;
            15'b11101011_1111_101: DATA = 1'b0;
            15'b11101011_1111_110: DATA = 1'b1;
            15'b11101011_1111_111: DATA = 1'b1;
            default: DATA = 1'b0;
        endcase
    end
endmodule
