`timescale 1ns / 1ps

module dds_sine_rom(
    input CLK,
    input [11:0] PHASE,
    input [1:0] FORM,
    output reg [11:0] DATA
    );
    
    reg [11:0] PHASE_REG;
    reg [1:0] FORM_REG;
    
    always @ (posedge CLK) begin
        PHASE_REG <= PHASE;
        FORM_REG <= FORM;
    end
    
    always @ (*) begin
        case ({FORM_REG, PHASE_REG})
            14'b00_000000000000: DATA = 12'b100000000000;
            14'b00_000000000001: DATA = 12'b100000000011;
            14'b00_000000000010: DATA = 12'b100000000110;
            14'b00_000000000011: DATA = 12'b100000001001;
            14'b00_000000000100: DATA = 12'b100000001100;
            14'b00_000000000101: DATA = 12'b100000001111;
            14'b00_000000000110: DATA = 12'b100000010010;
            14'b00_000000000111: DATA = 12'b100000010101;
            14'b00_000000001000: DATA = 12'b100000011001;
            14'b00_000000001001: DATA = 12'b100000011100;
            14'b00_000000001010: DATA = 12'b100000011111;
            14'b00_000000001011: DATA = 12'b100000100010;
            14'b00_000000001100: DATA = 12'b100000100101;
            14'b00_000000001101: DATA = 12'b100000101000;
            14'b00_000000001110: DATA = 12'b100000101011;
            14'b00_000000001111: DATA = 12'b100000101111;
            14'b00_000000010000: DATA = 12'b100000110010;
            14'b00_000000010001: DATA = 12'b100000110101;
            14'b00_000000010010: DATA = 12'b100000111000;
            14'b00_000000010011: DATA = 12'b100000111011;
            14'b00_000000010100: DATA = 12'b100000111110;
            14'b00_000000010101: DATA = 12'b100001000001;
            14'b00_000000010110: DATA = 12'b100001000101;
            14'b00_000000010111: DATA = 12'b100001001000;
            14'b00_000000011000: DATA = 12'b100001001011;
            14'b00_000000011001: DATA = 12'b100001001110;
            14'b00_000000011010: DATA = 12'b100001010001;
            14'b00_000000011011: DATA = 12'b100001010100;
            14'b00_000000011100: DATA = 12'b100001010111;
            14'b00_000000011101: DATA = 12'b100001011011;
            14'b00_000000011110: DATA = 12'b100001011110;
            14'b00_000000011111: DATA = 12'b100001100001;
            14'b00_000000100000: DATA = 12'b100001100100;
            14'b00_000000100001: DATA = 12'b100001100111;
            14'b00_000000100010: DATA = 12'b100001101010;
            14'b00_000000100011: DATA = 12'b100001101101;
            14'b00_000000100100: DATA = 12'b100001110000;
            14'b00_000000100101: DATA = 12'b100001110100;
            14'b00_000000100110: DATA = 12'b100001110111;
            14'b00_000000100111: DATA = 12'b100001111010;
            14'b00_000000101000: DATA = 12'b100001111101;
            14'b00_000000101001: DATA = 12'b100010000000;
            14'b00_000000101010: DATA = 12'b100010000011;
            14'b00_000000101011: DATA = 12'b100010000110;
            14'b00_000000101100: DATA = 12'b100010001010;
            14'b00_000000101101: DATA = 12'b100010001101;
            14'b00_000000101110: DATA = 12'b100010010000;
            14'b00_000000101111: DATA = 12'b100010010011;
            14'b00_000000110000: DATA = 12'b100010010110;
            14'b00_000000110001: DATA = 12'b100010011001;
            14'b00_000000110010: DATA = 12'b100010011100;
            14'b00_000000110011: DATA = 12'b100010011111;
            14'b00_000000110100: DATA = 12'b100010100011;
            14'b00_000000110101: DATA = 12'b100010100110;
            14'b00_000000110110: DATA = 12'b100010101001;
            14'b00_000000110111: DATA = 12'b100010101100;
            14'b00_000000111000: DATA = 12'b100010101111;
            14'b00_000000111001: DATA = 12'b100010110010;
            14'b00_000000111010: DATA = 12'b100010110101;
            14'b00_000000111011: DATA = 12'b100010111001;
            14'b00_000000111100: DATA = 12'b100010111100;
            14'b00_000000111101: DATA = 12'b100010111111;
            14'b00_000000111110: DATA = 12'b100011000010;
            14'b00_000000111111: DATA = 12'b100011000101;
            14'b00_000001000000: DATA = 12'b100011001000;
            14'b00_000001000001: DATA = 12'b100011001011;
            14'b00_000001000010: DATA = 12'b100011001110;
            14'b00_000001000011: DATA = 12'b100011010010;
            14'b00_000001000100: DATA = 12'b100011010101;
            14'b00_000001000101: DATA = 12'b100011011000;
            14'b00_000001000110: DATA = 12'b100011011011;
            14'b00_000001000111: DATA = 12'b100011011110;
            14'b00_000001001000: DATA = 12'b100011100001;
            14'b00_000001001001: DATA = 12'b100011100100;
            14'b00_000001001010: DATA = 12'b100011100111;
            14'b00_000001001011: DATA = 12'b100011101010;
            14'b00_000001001100: DATA = 12'b100011101110;
            14'b00_000001001101: DATA = 12'b100011110001;
            14'b00_000001001110: DATA = 12'b100011110100;
            14'b00_000001001111: DATA = 12'b100011110111;
            14'b00_000001010000: DATA = 12'b100011111010;
            14'b00_000001010001: DATA = 12'b100011111101;
            14'b00_000001010010: DATA = 12'b100100000000;
            14'b00_000001010011: DATA = 12'b100100000011;
            14'b00_000001010100: DATA = 12'b100100000111;
            14'b00_000001010101: DATA = 12'b100100001010;
            14'b00_000001010110: DATA = 12'b100100001101;
            14'b00_000001010111: DATA = 12'b100100010000;
            14'b00_000001011000: DATA = 12'b100100010011;
            14'b00_000001011001: DATA = 12'b100100010110;
            14'b00_000001011010: DATA = 12'b100100011001;
            14'b00_000001011011: DATA = 12'b100100011100;
            14'b00_000001011100: DATA = 12'b100100011111;
            14'b00_000001011101: DATA = 12'b100100100011;
            14'b00_000001011110: DATA = 12'b100100100110;
            14'b00_000001011111: DATA = 12'b100100101001;
            14'b00_000001100000: DATA = 12'b100100101100;
            14'b00_000001100001: DATA = 12'b100100101111;
            14'b00_000001100010: DATA = 12'b100100110010;
            14'b00_000001100011: DATA = 12'b100100110101;
            14'b00_000001100100: DATA = 12'b100100111000;
            14'b00_000001100101: DATA = 12'b100100111011;
            14'b00_000001100110: DATA = 12'b100100111110;
            14'b00_000001100111: DATA = 12'b100101000010;
            14'b00_000001101000: DATA = 12'b100101000101;
            14'b00_000001101001: DATA = 12'b100101001000;
            14'b00_000001101010: DATA = 12'b100101001011;
            14'b00_000001101011: DATA = 12'b100101001110;
            14'b00_000001101100: DATA = 12'b100101010001;
            14'b00_000001101101: DATA = 12'b100101010100;
            14'b00_000001101110: DATA = 12'b100101010111;
            14'b00_000001101111: DATA = 12'b100101011010;
            14'b00_000001110000: DATA = 12'b100101011101;
            14'b00_000001110001: DATA = 12'b100101100001;
            14'b00_000001110010: DATA = 12'b100101100100;
            14'b00_000001110011: DATA = 12'b100101100111;
            14'b00_000001110100: DATA = 12'b100101101010;
            14'b00_000001110101: DATA = 12'b100101101101;
            14'b00_000001110110: DATA = 12'b100101110000;
            14'b00_000001110111: DATA = 12'b100101110011;
            14'b00_000001111000: DATA = 12'b100101110110;
            14'b00_000001111001: DATA = 12'b100101111001;
            14'b00_000001111010: DATA = 12'b100101111100;
            14'b00_000001111011: DATA = 12'b100101111111;
            14'b00_000001111100: DATA = 12'b100110000011;
            14'b00_000001111101: DATA = 12'b100110000110;
            14'b00_000001111110: DATA = 12'b100110001001;
            14'b00_000001111111: DATA = 12'b100110001100;
            14'b00_000010000000: DATA = 12'b100110001111;
            14'b00_000010000001: DATA = 12'b100110010010;
            14'b00_000010000010: DATA = 12'b100110010101;
            14'b00_000010000011: DATA = 12'b100110011000;
            14'b00_000010000100: DATA = 12'b100110011011;
            14'b00_000010000101: DATA = 12'b100110011110;
            14'b00_000010000110: DATA = 12'b100110100001;
            14'b00_000010000111: DATA = 12'b100110100100;
            14'b00_000010001000: DATA = 12'b100110100111;
            14'b00_000010001001: DATA = 12'b100110101011;
            14'b00_000010001010: DATA = 12'b100110101110;
            14'b00_000010001011: DATA = 12'b100110110001;
            14'b00_000010001100: DATA = 12'b100110110100;
            14'b00_000010001101: DATA = 12'b100110110111;
            14'b00_000010001110: DATA = 12'b100110111010;
            14'b00_000010001111: DATA = 12'b100110111101;
            14'b00_000010010000: DATA = 12'b100111000000;
            14'b00_000010010001: DATA = 12'b100111000011;
            14'b00_000010010010: DATA = 12'b100111000110;
            14'b00_000010010011: DATA = 12'b100111001001;
            14'b00_000010010100: DATA = 12'b100111001100;
            14'b00_000010010101: DATA = 12'b100111001111;
            14'b00_000010010110: DATA = 12'b100111010010;
            14'b00_000010010111: DATA = 12'b100111010101;
            14'b00_000010011000: DATA = 12'b100111011000;
            14'b00_000010011001: DATA = 12'b100111011100;
            14'b00_000010011010: DATA = 12'b100111011111;
            14'b00_000010011011: DATA = 12'b100111100010;
            14'b00_000010011100: DATA = 12'b100111100101;
            14'b00_000010011101: DATA = 12'b100111101000;
            14'b00_000010011110: DATA = 12'b100111101011;
            14'b00_000010011111: DATA = 12'b100111101110;
            14'b00_000010100000: DATA = 12'b100111110001;
            14'b00_000010100001: DATA = 12'b100111110100;
            14'b00_000010100010: DATA = 12'b100111110111;
            14'b00_000010100011: DATA = 12'b100111111010;
            14'b00_000010100100: DATA = 12'b100111111101;
            14'b00_000010100101: DATA = 12'b101000000000;
            14'b00_000010100110: DATA = 12'b101000000011;
            14'b00_000010100111: DATA = 12'b101000000110;
            14'b00_000010101000: DATA = 12'b101000001001;
            14'b00_000010101001: DATA = 12'b101000001100;
            14'b00_000010101010: DATA = 12'b101000001111;
            14'b00_000010101011: DATA = 12'b101000010010;
            14'b00_000010101100: DATA = 12'b101000010101;
            14'b00_000010101101: DATA = 12'b101000011000;
            14'b00_000010101110: DATA = 12'b101000011011;
            14'b00_000010101111: DATA = 12'b101000011110;
            14'b00_000010110000: DATA = 12'b101000100001;
            14'b00_000010110001: DATA = 12'b101000100100;
            14'b00_000010110010: DATA = 12'b101000101000;
            14'b00_000010110011: DATA = 12'b101000101011;
            14'b00_000010110100: DATA = 12'b101000101110;
            14'b00_000010110101: DATA = 12'b101000110001;
            14'b00_000010110110: DATA = 12'b101000110100;
            14'b00_000010110111: DATA = 12'b101000110111;
            14'b00_000010111000: DATA = 12'b101000111010;
            14'b00_000010111001: DATA = 12'b101000111101;
            14'b00_000010111010: DATA = 12'b101001000000;
            14'b00_000010111011: DATA = 12'b101001000011;
            14'b00_000010111100: DATA = 12'b101001000110;
            14'b00_000010111101: DATA = 12'b101001001001;
            14'b00_000010111110: DATA = 12'b101001001100;
            14'b00_000010111111: DATA = 12'b101001001111;
            14'b00_000011000000: DATA = 12'b101001010010;
            14'b00_000011000001: DATA = 12'b101001010101;
            14'b00_000011000010: DATA = 12'b101001011000;
            14'b00_000011000011: DATA = 12'b101001011011;
            14'b00_000011000100: DATA = 12'b101001011110;
            14'b00_000011000101: DATA = 12'b101001100001;
            14'b00_000011000110: DATA = 12'b101001100100;
            14'b00_000011000111: DATA = 12'b101001100111;
            14'b00_000011001000: DATA = 12'b101001101010;
            14'b00_000011001001: DATA = 12'b101001101101;
            14'b00_000011001010: DATA = 12'b101001110000;
            14'b00_000011001011: DATA = 12'b101001110011;
            14'b00_000011001100: DATA = 12'b101001110110;
            14'b00_000011001101: DATA = 12'b101001111001;
            14'b00_000011001110: DATA = 12'b101001111100;
            14'b00_000011001111: DATA = 12'b101001111111;
            14'b00_000011010000: DATA = 12'b101010000010;
            14'b00_000011010001: DATA = 12'b101010000101;
            14'b00_000011010010: DATA = 12'b101010001000;
            14'b00_000011010011: DATA = 12'b101010001011;
            14'b00_000011010100: DATA = 12'b101010001110;
            14'b00_000011010101: DATA = 12'b101010010000;
            14'b00_000011010110: DATA = 12'b101010010011;
            14'b00_000011010111: DATA = 12'b101010010110;
            14'b00_000011011000: DATA = 12'b101010011001;
            14'b00_000011011001: DATA = 12'b101010011100;
            14'b00_000011011010: DATA = 12'b101010011111;
            14'b00_000011011011: DATA = 12'b101010100010;
            14'b00_000011011100: DATA = 12'b101010100101;
            14'b00_000011011101: DATA = 12'b101010101000;
            14'b00_000011011110: DATA = 12'b101010101011;
            14'b00_000011011111: DATA = 12'b101010101110;
            14'b00_000011100000: DATA = 12'b101010110001;
            14'b00_000011100001: DATA = 12'b101010110100;
            14'b00_000011100010: DATA = 12'b101010110111;
            14'b00_000011100011: DATA = 12'b101010111010;
            14'b00_000011100100: DATA = 12'b101010111101;
            14'b00_000011100101: DATA = 12'b101011000000;
            14'b00_000011100110: DATA = 12'b101011000011;
            14'b00_000011100111: DATA = 12'b101011000110;
            14'b00_000011101000: DATA = 12'b101011001001;
            14'b00_000011101001: DATA = 12'b101011001100;
            14'b00_000011101010: DATA = 12'b101011001111;
            14'b00_000011101011: DATA = 12'b101011010010;
            14'b00_000011101100: DATA = 12'b101011010100;
            14'b00_000011101101: DATA = 12'b101011010111;
            14'b00_000011101110: DATA = 12'b101011011010;
            14'b00_000011101111: DATA = 12'b101011011101;
            14'b00_000011110000: DATA = 12'b101011100000;
            14'b00_000011110001: DATA = 12'b101011100011;
            14'b00_000011110010: DATA = 12'b101011100110;
            14'b00_000011110011: DATA = 12'b101011101001;
            14'b00_000011110100: DATA = 12'b101011101100;
            14'b00_000011110101: DATA = 12'b101011101111;
            14'b00_000011110110: DATA = 12'b101011110010;
            14'b00_000011110111: DATA = 12'b101011110101;
            14'b00_000011111000: DATA = 12'b101011111000;
            14'b00_000011111001: DATA = 12'b101011111011;
            14'b00_000011111010: DATA = 12'b101011111101;
            14'b00_000011111011: DATA = 12'b101100000000;
            14'b00_000011111100: DATA = 12'b101100000011;
            14'b00_000011111101: DATA = 12'b101100000110;
            14'b00_000011111110: DATA = 12'b101100001001;
            14'b00_000011111111: DATA = 12'b101100001100;
            14'b00_000100000000: DATA = 12'b101100001111;
            14'b00_000100000001: DATA = 12'b101100010010;
            14'b00_000100000010: DATA = 12'b101100010101;
            14'b00_000100000011: DATA = 12'b101100011000;
            14'b00_000100000100: DATA = 12'b101100011010;
            14'b00_000100000101: DATA = 12'b101100011101;
            14'b00_000100000110: DATA = 12'b101100100000;
            14'b00_000100000111: DATA = 12'b101100100011;
            14'b00_000100001000: DATA = 12'b101100100110;
            14'b00_000100001001: DATA = 12'b101100101001;
            14'b00_000100001010: DATA = 12'b101100101100;
            14'b00_000100001011: DATA = 12'b101100101111;
            14'b00_000100001100: DATA = 12'b101100110010;
            14'b00_000100001101: DATA = 12'b101100110100;
            14'b00_000100001110: DATA = 12'b101100110111;
            14'b00_000100001111: DATA = 12'b101100111010;
            14'b00_000100010000: DATA = 12'b101100111101;
            14'b00_000100010001: DATA = 12'b101101000000;
            14'b00_000100010010: DATA = 12'b101101000011;
            14'b00_000100010011: DATA = 12'b101101000110;
            14'b00_000100010100: DATA = 12'b101101001000;
            14'b00_000100010101: DATA = 12'b101101001011;
            14'b00_000100010110: DATA = 12'b101101001110;
            14'b00_000100010111: DATA = 12'b101101010001;
            14'b00_000100011000: DATA = 12'b101101010100;
            14'b00_000100011001: DATA = 12'b101101010111;
            14'b00_000100011010: DATA = 12'b101101011010;
            14'b00_000100011011: DATA = 12'b101101011100;
            14'b00_000100011100: DATA = 12'b101101011111;
            14'b00_000100011101: DATA = 12'b101101100010;
            14'b00_000100011110: DATA = 12'b101101100101;
            14'b00_000100011111: DATA = 12'b101101101000;
            14'b00_000100100000: DATA = 12'b101101101011;
            14'b00_000100100001: DATA = 12'b101101101110;
            14'b00_000100100010: DATA = 12'b101101110000;
            14'b00_000100100011: DATA = 12'b101101110011;
            14'b00_000100100100: DATA = 12'b101101110110;
            14'b00_000100100101: DATA = 12'b101101111001;
            14'b00_000100100110: DATA = 12'b101101111100;
            14'b00_000100100111: DATA = 12'b101101111111;
            14'b00_000100101000: DATA = 12'b101110000001;
            14'b00_000100101001: DATA = 12'b101110000100;
            14'b00_000100101010: DATA = 12'b101110000111;
            14'b00_000100101011: DATA = 12'b101110001010;
            14'b00_000100101100: DATA = 12'b101110001101;
            14'b00_000100101101: DATA = 12'b101110001111;
            14'b00_000100101110: DATA = 12'b101110010010;
            14'b00_000100101111: DATA = 12'b101110010101;
            14'b00_000100110000: DATA = 12'b101110011000;
            14'b00_000100110001: DATA = 12'b101110011011;
            14'b00_000100110010: DATA = 12'b101110011101;
            14'b00_000100110011: DATA = 12'b101110100000;
            14'b00_000100110100: DATA = 12'b101110100011;
            14'b00_000100110101: DATA = 12'b101110100110;
            14'b00_000100110110: DATA = 12'b101110101001;
            14'b00_000100110111: DATA = 12'b101110101011;
            14'b00_000100111000: DATA = 12'b101110101110;
            14'b00_000100111001: DATA = 12'b101110110001;
            14'b00_000100111010: DATA = 12'b101110110100;
            14'b00_000100111011: DATA = 12'b101110110111;
            14'b00_000100111100: DATA = 12'b101110111001;
            14'b00_000100111101: DATA = 12'b101110111100;
            14'b00_000100111110: DATA = 12'b101110111111;
            14'b00_000100111111: DATA = 12'b101111000010;
            14'b00_000101000000: DATA = 12'b101111000100;
            14'b00_000101000001: DATA = 12'b101111000111;
            14'b00_000101000010: DATA = 12'b101111001010;
            14'b00_000101000011: DATA = 12'b101111001101;
            14'b00_000101000100: DATA = 12'b101111010000;
            14'b00_000101000101: DATA = 12'b101111010010;
            14'b00_000101000110: DATA = 12'b101111010101;
            14'b00_000101000111: DATA = 12'b101111011000;
            14'b00_000101001000: DATA = 12'b101111011011;
            14'b00_000101001001: DATA = 12'b101111011101;
            14'b00_000101001010: DATA = 12'b101111100000;
            14'b00_000101001011: DATA = 12'b101111100011;
            14'b00_000101001100: DATA = 12'b101111100110;
            14'b00_000101001101: DATA = 12'b101111101000;
            14'b00_000101001110: DATA = 12'b101111101011;
            14'b00_000101001111: DATA = 12'b101111101110;
            14'b00_000101010000: DATA = 12'b101111110000;
            14'b00_000101010001: DATA = 12'b101111110011;
            14'b00_000101010010: DATA = 12'b101111110110;
            14'b00_000101010011: DATA = 12'b101111111001;
            14'b00_000101010100: DATA = 12'b101111111011;
            14'b00_000101010101: DATA = 12'b101111111110;
            14'b00_000101010110: DATA = 12'b110000000001;
            14'b00_000101010111: DATA = 12'b110000000100;
            14'b00_000101011000: DATA = 12'b110000000110;
            14'b00_000101011001: DATA = 12'b110000001001;
            14'b00_000101011010: DATA = 12'b110000001100;
            14'b00_000101011011: DATA = 12'b110000001110;
            14'b00_000101011100: DATA = 12'b110000010001;
            14'b00_000101011101: DATA = 12'b110000010100;
            14'b00_000101011110: DATA = 12'b110000010110;
            14'b00_000101011111: DATA = 12'b110000011001;
            14'b00_000101100000: DATA = 12'b110000011100;
            14'b00_000101100001: DATA = 12'b110000011111;
            14'b00_000101100010: DATA = 12'b110000100001;
            14'b00_000101100011: DATA = 12'b110000100100;
            14'b00_000101100100: DATA = 12'b110000100111;
            14'b00_000101100101: DATA = 12'b110000101001;
            14'b00_000101100110: DATA = 12'b110000101100;
            14'b00_000101100111: DATA = 12'b110000101111;
            14'b00_000101101000: DATA = 12'b110000110001;
            14'b00_000101101001: DATA = 12'b110000110100;
            14'b00_000101101010: DATA = 12'b110000110111;
            14'b00_000101101011: DATA = 12'b110000111001;
            14'b00_000101101100: DATA = 12'b110000111100;
            14'b00_000101101101: DATA = 12'b110000111111;
            14'b00_000101101110: DATA = 12'b110001000001;
            14'b00_000101101111: DATA = 12'b110001000100;
            14'b00_000101110000: DATA = 12'b110001000111;
            14'b00_000101110001: DATA = 12'b110001001001;
            14'b00_000101110010: DATA = 12'b110001001100;
            14'b00_000101110011: DATA = 12'b110001001111;
            14'b00_000101110100: DATA = 12'b110001010001;
            14'b00_000101110101: DATA = 12'b110001010100;
            14'b00_000101110110: DATA = 12'b110001010111;
            14'b00_000101110111: DATA = 12'b110001011001;
            14'b00_000101111000: DATA = 12'b110001011100;
            14'b00_000101111001: DATA = 12'b110001011110;
            14'b00_000101111010: DATA = 12'b110001100001;
            14'b00_000101111011: DATA = 12'b110001100100;
            14'b00_000101111100: DATA = 12'b110001100110;
            14'b00_000101111101: DATA = 12'b110001101001;
            14'b00_000101111110: DATA = 12'b110001101100;
            14'b00_000101111111: DATA = 12'b110001101110;
            14'b00_000110000000: DATA = 12'b110001110001;
            14'b00_000110000001: DATA = 12'b110001110011;
            14'b00_000110000010: DATA = 12'b110001110110;
            14'b00_000110000011: DATA = 12'b110001111001;
            14'b00_000110000100: DATA = 12'b110001111011;
            14'b00_000110000101: DATA = 12'b110001111110;
            14'b00_000110000110: DATA = 12'b110010000000;
            14'b00_000110000111: DATA = 12'b110010000011;
            14'b00_000110001000: DATA = 12'b110010000110;
            14'b00_000110001001: DATA = 12'b110010001000;
            14'b00_000110001010: DATA = 12'b110010001011;
            14'b00_000110001011: DATA = 12'b110010001101;
            14'b00_000110001100: DATA = 12'b110010010000;
            14'b00_000110001101: DATA = 12'b110010010010;
            14'b00_000110001110: DATA = 12'b110010010101;
            14'b00_000110001111: DATA = 12'b110010011000;
            14'b00_000110010000: DATA = 12'b110010011010;
            14'b00_000110010001: DATA = 12'b110010011101;
            14'b00_000110010010: DATA = 12'b110010011111;
            14'b00_000110010011: DATA = 12'b110010100010;
            14'b00_000110010100: DATA = 12'b110010100100;
            14'b00_000110010101: DATA = 12'b110010100111;
            14'b00_000110010110: DATA = 12'b110010101010;
            14'b00_000110010111: DATA = 12'b110010101100;
            14'b00_000110011000: DATA = 12'b110010101111;
            14'b00_000110011001: DATA = 12'b110010110001;
            14'b00_000110011010: DATA = 12'b110010110100;
            14'b00_000110011011: DATA = 12'b110010110110;
            14'b00_000110011100: DATA = 12'b110010111001;
            14'b00_000110011101: DATA = 12'b110010111011;
            14'b00_000110011110: DATA = 12'b110010111110;
            14'b00_000110011111: DATA = 12'b110011000000;
            14'b00_000110100000: DATA = 12'b110011000011;
            14'b00_000110100001: DATA = 12'b110011000101;
            14'b00_000110100010: DATA = 12'b110011001000;
            14'b00_000110100011: DATA = 12'b110011001010;
            14'b00_000110100100: DATA = 12'b110011001101;
            14'b00_000110100101: DATA = 12'b110011001111;
            14'b00_000110100110: DATA = 12'b110011010010;
            14'b00_000110100111: DATA = 12'b110011010100;
            14'b00_000110101000: DATA = 12'b110011010111;
            14'b00_000110101001: DATA = 12'b110011011001;
            14'b00_000110101010: DATA = 12'b110011011100;
            14'b00_000110101011: DATA = 12'b110011011110;
            14'b00_000110101100: DATA = 12'b110011100001;
            14'b00_000110101101: DATA = 12'b110011100011;
            14'b00_000110101110: DATA = 12'b110011100110;
            14'b00_000110101111: DATA = 12'b110011101000;
            14'b00_000110110000: DATA = 12'b110011101011;
            14'b00_000110110001: DATA = 12'b110011101101;
            14'b00_000110110010: DATA = 12'b110011110000;
            14'b00_000110110011: DATA = 12'b110011110010;
            14'b00_000110110100: DATA = 12'b110011110101;
            14'b00_000110110101: DATA = 12'b110011110111;
            14'b00_000110110110: DATA = 12'b110011111010;
            14'b00_000110110111: DATA = 12'b110011111100;
            14'b00_000110111000: DATA = 12'b110011111111;
            14'b00_000110111001: DATA = 12'b110100000001;
            14'b00_000110111010: DATA = 12'b110100000011;
            14'b00_000110111011: DATA = 12'b110100000110;
            14'b00_000110111100: DATA = 12'b110100001000;
            14'b00_000110111101: DATA = 12'b110100001011;
            14'b00_000110111110: DATA = 12'b110100001101;
            14'b00_000110111111: DATA = 12'b110100010000;
            14'b00_000111000000: DATA = 12'b110100010010;
            14'b00_000111000001: DATA = 12'b110100010101;
            14'b00_000111000010: DATA = 12'b110100010111;
            14'b00_000111000011: DATA = 12'b110100011001;
            14'b00_000111000100: DATA = 12'b110100011100;
            14'b00_000111000101: DATA = 12'b110100011110;
            14'b00_000111000110: DATA = 12'b110100100001;
            14'b00_000111000111: DATA = 12'b110100100011;
            14'b00_000111001000: DATA = 12'b110100100101;
            14'b00_000111001001: DATA = 12'b110100101000;
            14'b00_000111001010: DATA = 12'b110100101010;
            14'b00_000111001011: DATA = 12'b110100101101;
            14'b00_000111001100: DATA = 12'b110100101111;
            14'b00_000111001101: DATA = 12'b110100110001;
            14'b00_000111001110: DATA = 12'b110100110100;
            14'b00_000111001111: DATA = 12'b110100110110;
            14'b00_000111010000: DATA = 12'b110100111001;
            14'b00_000111010001: DATA = 12'b110100111011;
            14'b00_000111010010: DATA = 12'b110100111101;
            14'b00_000111010011: DATA = 12'b110101000000;
            14'b00_000111010100: DATA = 12'b110101000010;
            14'b00_000111010101: DATA = 12'b110101000100;
            14'b00_000111010110: DATA = 12'b110101000111;
            14'b00_000111010111: DATA = 12'b110101001001;
            14'b00_000111011000: DATA = 12'b110101001011;
            14'b00_000111011001: DATA = 12'b110101001110;
            14'b00_000111011010: DATA = 12'b110101010000;
            14'b00_000111011011: DATA = 12'b110101010011;
            14'b00_000111011100: DATA = 12'b110101010101;
            14'b00_000111011101: DATA = 12'b110101010111;
            14'b00_000111011110: DATA = 12'b110101011010;
            14'b00_000111011111: DATA = 12'b110101011100;
            14'b00_000111100000: DATA = 12'b110101011110;
            14'b00_000111100001: DATA = 12'b110101100001;
            14'b00_000111100010: DATA = 12'b110101100011;
            14'b00_000111100011: DATA = 12'b110101100101;
            14'b00_000111100100: DATA = 12'b110101100111;
            14'b00_000111100101: DATA = 12'b110101101010;
            14'b00_000111100110: DATA = 12'b110101101100;
            14'b00_000111100111: DATA = 12'b110101101110;
            14'b00_000111101000: DATA = 12'b110101110001;
            14'b00_000111101001: DATA = 12'b110101110011;
            14'b00_000111101010: DATA = 12'b110101110101;
            14'b00_000111101011: DATA = 12'b110101111000;
            14'b00_000111101100: DATA = 12'b110101111010;
            14'b00_000111101101: DATA = 12'b110101111100;
            14'b00_000111101110: DATA = 12'b110101111110;
            14'b00_000111101111: DATA = 12'b110110000001;
            14'b00_000111110000: DATA = 12'b110110000011;
            14'b00_000111110001: DATA = 12'b110110000101;
            14'b00_000111110010: DATA = 12'b110110001000;
            14'b00_000111110011: DATA = 12'b110110001010;
            14'b00_000111110100: DATA = 12'b110110001100;
            14'b00_000111110101: DATA = 12'b110110001110;
            14'b00_000111110110: DATA = 12'b110110010001;
            14'b00_000111110111: DATA = 12'b110110010011;
            14'b00_000111111000: DATA = 12'b110110010101;
            14'b00_000111111001: DATA = 12'b110110010111;
            14'b00_000111111010: DATA = 12'b110110011010;
            14'b00_000111111011: DATA = 12'b110110011100;
            14'b00_000111111100: DATA = 12'b110110011110;
            14'b00_000111111101: DATA = 12'b110110100000;
            14'b00_000111111110: DATA = 12'b110110100011;
            14'b00_000111111111: DATA = 12'b110110100101;
            14'b00_001000000000: DATA = 12'b110110100111;
            14'b00_001000000001: DATA = 12'b110110101001;
            14'b00_001000000010: DATA = 12'b110110101011;
            14'b00_001000000011: DATA = 12'b110110101110;
            14'b00_001000000100: DATA = 12'b110110110000;
            14'b00_001000000101: DATA = 12'b110110110010;
            14'b00_001000000110: DATA = 12'b110110110100;
            14'b00_001000000111: DATA = 12'b110110110110;
            14'b00_001000001000: DATA = 12'b110110111001;
            14'b00_001000001001: DATA = 12'b110110111011;
            14'b00_001000001010: DATA = 12'b110110111101;
            14'b00_001000001011: DATA = 12'b110110111111;
            14'b00_001000001100: DATA = 12'b110111000001;
            14'b00_001000001101: DATA = 12'b110111000100;
            14'b00_001000001110: DATA = 12'b110111000110;
            14'b00_001000001111: DATA = 12'b110111001000;
            14'b00_001000010000: DATA = 12'b110111001010;
            14'b00_001000010001: DATA = 12'b110111001100;
            14'b00_001000010010: DATA = 12'b110111001110;
            14'b00_001000010011: DATA = 12'b110111010001;
            14'b00_001000010100: DATA = 12'b110111010011;
            14'b00_001000010101: DATA = 12'b110111010101;
            14'b00_001000010110: DATA = 12'b110111010111;
            14'b00_001000010111: DATA = 12'b110111011001;
            14'b00_001000011000: DATA = 12'b110111011011;
            14'b00_001000011001: DATA = 12'b110111011101;
            14'b00_001000011010: DATA = 12'b110111100000;
            14'b00_001000011011: DATA = 12'b110111100010;
            14'b00_001000011100: DATA = 12'b110111100100;
            14'b00_001000011101: DATA = 12'b110111100110;
            14'b00_001000011110: DATA = 12'b110111101000;
            14'b00_001000011111: DATA = 12'b110111101010;
            14'b00_001000100000: DATA = 12'b110111101100;
            14'b00_001000100001: DATA = 12'b110111101110;
            14'b00_001000100010: DATA = 12'b110111110000;
            14'b00_001000100011: DATA = 12'b110111110011;
            14'b00_001000100100: DATA = 12'b110111110101;
            14'b00_001000100101: DATA = 12'b110111110111;
            14'b00_001000100110: DATA = 12'b110111111001;
            14'b00_001000100111: DATA = 12'b110111111011;
            14'b00_001000101000: DATA = 12'b110111111101;
            14'b00_001000101001: DATA = 12'b110111111111;
            14'b00_001000101010: DATA = 12'b111000000001;
            14'b00_001000101011: DATA = 12'b111000000011;
            14'b00_001000101100: DATA = 12'b111000000101;
            14'b00_001000101101: DATA = 12'b111000000111;
            14'b00_001000101110: DATA = 12'b111000001001;
            14'b00_001000101111: DATA = 12'b111000001011;
            14'b00_001000110000: DATA = 12'b111000001110;
            14'b00_001000110001: DATA = 12'b111000010000;
            14'b00_001000110010: DATA = 12'b111000010010;
            14'b00_001000110011: DATA = 12'b111000010100;
            14'b00_001000110100: DATA = 12'b111000010110;
            14'b00_001000110101: DATA = 12'b111000011000;
            14'b00_001000110110: DATA = 12'b111000011010;
            14'b00_001000110111: DATA = 12'b111000011100;
            14'b00_001000111000: DATA = 12'b111000011110;
            14'b00_001000111001: DATA = 12'b111000100000;
            14'b00_001000111010: DATA = 12'b111000100010;
            14'b00_001000111011: DATA = 12'b111000100100;
            14'b00_001000111100: DATA = 12'b111000100110;
            14'b00_001000111101: DATA = 12'b111000101000;
            14'b00_001000111110: DATA = 12'b111000101010;
            14'b00_001000111111: DATA = 12'b111000101100;
            14'b00_001001000000: DATA = 12'b111000101110;
            14'b00_001001000001: DATA = 12'b111000110000;
            14'b00_001001000010: DATA = 12'b111000110010;
            14'b00_001001000011: DATA = 12'b111000110100;
            14'b00_001001000100: DATA = 12'b111000110110;
            14'b00_001001000101: DATA = 12'b111000111000;
            14'b00_001001000110: DATA = 12'b111000111010;
            14'b00_001001000111: DATA = 12'b111000111100;
            14'b00_001001001000: DATA = 12'b111000111110;
            14'b00_001001001001: DATA = 12'b111001000000;
            14'b00_001001001010: DATA = 12'b111001000010;
            14'b00_001001001011: DATA = 12'b111001000100;
            14'b00_001001001100: DATA = 12'b111001000101;
            14'b00_001001001101: DATA = 12'b111001000111;
            14'b00_001001001110: DATA = 12'b111001001001;
            14'b00_001001001111: DATA = 12'b111001001011;
            14'b00_001001010000: DATA = 12'b111001001101;
            14'b00_001001010001: DATA = 12'b111001001111;
            14'b00_001001010010: DATA = 12'b111001010001;
            14'b00_001001010011: DATA = 12'b111001010011;
            14'b00_001001010100: DATA = 12'b111001010101;
            14'b00_001001010101: DATA = 12'b111001010111;
            14'b00_001001010110: DATA = 12'b111001011001;
            14'b00_001001010111: DATA = 12'b111001011011;
            14'b00_001001011000: DATA = 12'b111001011101;
            14'b00_001001011001: DATA = 12'b111001011110;
            14'b00_001001011010: DATA = 12'b111001100000;
            14'b00_001001011011: DATA = 12'b111001100010;
            14'b00_001001011100: DATA = 12'b111001100100;
            14'b00_001001011101: DATA = 12'b111001100110;
            14'b00_001001011110: DATA = 12'b111001101000;
            14'b00_001001011111: DATA = 12'b111001101010;
            14'b00_001001100000: DATA = 12'b111001101100;
            14'b00_001001100001: DATA = 12'b111001101110;
            14'b00_001001100010: DATA = 12'b111001101111;
            14'b00_001001100011: DATA = 12'b111001110001;
            14'b00_001001100100: DATA = 12'b111001110011;
            14'b00_001001100101: DATA = 12'b111001110101;
            14'b00_001001100110: DATA = 12'b111001110111;
            14'b00_001001100111: DATA = 12'b111001111001;
            14'b00_001001101000: DATA = 12'b111001111011;
            14'b00_001001101001: DATA = 12'b111001111100;
            14'b00_001001101010: DATA = 12'b111001111110;
            14'b00_001001101011: DATA = 12'b111010000000;
            14'b00_001001101100: DATA = 12'b111010000010;
            14'b00_001001101101: DATA = 12'b111010000100;
            14'b00_001001101110: DATA = 12'b111010000101;
            14'b00_001001101111: DATA = 12'b111010000111;
            14'b00_001001110000: DATA = 12'b111010001001;
            14'b00_001001110001: DATA = 12'b111010001011;
            14'b00_001001110010: DATA = 12'b111010001101;
            14'b00_001001110011: DATA = 12'b111010001111;
            14'b00_001001110100: DATA = 12'b111010010000;
            14'b00_001001110101: DATA = 12'b111010010010;
            14'b00_001001110110: DATA = 12'b111010010100;
            14'b00_001001110111: DATA = 12'b111010010110;
            14'b00_001001111000: DATA = 12'b111010010111;
            14'b00_001001111001: DATA = 12'b111010011001;
            14'b00_001001111010: DATA = 12'b111010011011;
            14'b00_001001111011: DATA = 12'b111010011101;
            14'b00_001001111100: DATA = 12'b111010011111;
            14'b00_001001111101: DATA = 12'b111010100000;
            14'b00_001001111110: DATA = 12'b111010100010;
            14'b00_001001111111: DATA = 12'b111010100100;
            14'b00_001010000000: DATA = 12'b111010100110;
            14'b00_001010000001: DATA = 12'b111010100111;
            14'b00_001010000010: DATA = 12'b111010101001;
            14'b00_001010000011: DATA = 12'b111010101011;
            14'b00_001010000100: DATA = 12'b111010101100;
            14'b00_001010000101: DATA = 12'b111010101110;
            14'b00_001010000110: DATA = 12'b111010110000;
            14'b00_001010000111: DATA = 12'b111010110010;
            14'b00_001010001000: DATA = 12'b111010110011;
            14'b00_001010001001: DATA = 12'b111010110101;
            14'b00_001010001010: DATA = 12'b111010110111;
            14'b00_001010001011: DATA = 12'b111010111000;
            14'b00_001010001100: DATA = 12'b111010111010;
            14'b00_001010001101: DATA = 12'b111010111100;
            14'b00_001010001110: DATA = 12'b111010111110;
            14'b00_001010001111: DATA = 12'b111010111111;
            14'b00_001010010000: DATA = 12'b111011000001;
            14'b00_001010010001: DATA = 12'b111011000011;
            14'b00_001010010010: DATA = 12'b111011000100;
            14'b00_001010010011: DATA = 12'b111011000110;
            14'b00_001010010100: DATA = 12'b111011001000;
            14'b00_001010010101: DATA = 12'b111011001001;
            14'b00_001010010110: DATA = 12'b111011001011;
            14'b00_001010010111: DATA = 12'b111011001101;
            14'b00_001010011000: DATA = 12'b111011001110;
            14'b00_001010011001: DATA = 12'b111011010000;
            14'b00_001010011010: DATA = 12'b111011010010;
            14'b00_001010011011: DATA = 12'b111011010011;
            14'b00_001010011100: DATA = 12'b111011010101;
            14'b00_001010011101: DATA = 12'b111011010110;
            14'b00_001010011110: DATA = 12'b111011011000;
            14'b00_001010011111: DATA = 12'b111011011010;
            14'b00_001010100000: DATA = 12'b111011011011;
            14'b00_001010100001: DATA = 12'b111011011101;
            14'b00_001010100010: DATA = 12'b111011011110;
            14'b00_001010100011: DATA = 12'b111011100000;
            14'b00_001010100100: DATA = 12'b111011100010;
            14'b00_001010100101: DATA = 12'b111011100011;
            14'b00_001010100110: DATA = 12'b111011100101;
            14'b00_001010100111: DATA = 12'b111011100110;
            14'b00_001010101000: DATA = 12'b111011101000;
            14'b00_001010101001: DATA = 12'b111011101010;
            14'b00_001010101010: DATA = 12'b111011101011;
            14'b00_001010101011: DATA = 12'b111011101101;
            14'b00_001010101100: DATA = 12'b111011101110;
            14'b00_001010101101: DATA = 12'b111011110000;
            14'b00_001010101110: DATA = 12'b111011110001;
            14'b00_001010101111: DATA = 12'b111011110011;
            14'b00_001010110000: DATA = 12'b111011110101;
            14'b00_001010110001: DATA = 12'b111011110110;
            14'b00_001010110010: DATA = 12'b111011111000;
            14'b00_001010110011: DATA = 12'b111011111001;
            14'b00_001010110100: DATA = 12'b111011111011;
            14'b00_001010110101: DATA = 12'b111011111100;
            14'b00_001010110110: DATA = 12'b111011111110;
            14'b00_001010110111: DATA = 12'b111011111111;
            14'b00_001010111000: DATA = 12'b111100000001;
            14'b00_001010111001: DATA = 12'b111100000010;
            14'b00_001010111010: DATA = 12'b111100000100;
            14'b00_001010111011: DATA = 12'b111100000101;
            14'b00_001010111100: DATA = 12'b111100000111;
            14'b00_001010111101: DATA = 12'b111100001000;
            14'b00_001010111110: DATA = 12'b111100001010;
            14'b00_001010111111: DATA = 12'b111100001011;
            14'b00_001011000000: DATA = 12'b111100001101;
            14'b00_001011000001: DATA = 12'b111100001110;
            14'b00_001011000010: DATA = 12'b111100010000;
            14'b00_001011000011: DATA = 12'b111100010001;
            14'b00_001011000100: DATA = 12'b111100010011;
            14'b00_001011000101: DATA = 12'b111100010100;
            14'b00_001011000110: DATA = 12'b111100010110;
            14'b00_001011000111: DATA = 12'b111100010111;
            14'b00_001011001000: DATA = 12'b111100011000;
            14'b00_001011001001: DATA = 12'b111100011010;
            14'b00_001011001010: DATA = 12'b111100011011;
            14'b00_001011001011: DATA = 12'b111100011101;
            14'b00_001011001100: DATA = 12'b111100011110;
            14'b00_001011001101: DATA = 12'b111100100000;
            14'b00_001011001110: DATA = 12'b111100100001;
            14'b00_001011001111: DATA = 12'b111100100011;
            14'b00_001011010000: DATA = 12'b111100100100;
            14'b00_001011010001: DATA = 12'b111100100101;
            14'b00_001011010010: DATA = 12'b111100100111;
            14'b00_001011010011: DATA = 12'b111100101000;
            14'b00_001011010100: DATA = 12'b111100101010;
            14'b00_001011010101: DATA = 12'b111100101011;
            14'b00_001011010110: DATA = 12'b111100101100;
            14'b00_001011010111: DATA = 12'b111100101110;
            14'b00_001011011000: DATA = 12'b111100101111;
            14'b00_001011011001: DATA = 12'b111100110000;
            14'b00_001011011010: DATA = 12'b111100110010;
            14'b00_001011011011: DATA = 12'b111100110011;
            14'b00_001011011100: DATA = 12'b111100110101;
            14'b00_001011011101: DATA = 12'b111100110110;
            14'b00_001011011110: DATA = 12'b111100110111;
            14'b00_001011011111: DATA = 12'b111100111001;
            14'b00_001011100000: DATA = 12'b111100111010;
            14'b00_001011100001: DATA = 12'b111100111011;
            14'b00_001011100010: DATA = 12'b111100111101;
            14'b00_001011100011: DATA = 12'b111100111110;
            14'b00_001011100100: DATA = 12'b111100111111;
            14'b00_001011100101: DATA = 12'b111101000001;
            14'b00_001011100110: DATA = 12'b111101000010;
            14'b00_001011100111: DATA = 12'b111101000011;
            14'b00_001011101000: DATA = 12'b111101000101;
            14'b00_001011101001: DATA = 12'b111101000110;
            14'b00_001011101010: DATA = 12'b111101000111;
            14'b00_001011101011: DATA = 12'b111101001000;
            14'b00_001011101100: DATA = 12'b111101001010;
            14'b00_001011101101: DATA = 12'b111101001011;
            14'b00_001011101110: DATA = 12'b111101001100;
            14'b00_001011101111: DATA = 12'b111101001110;
            14'b00_001011110000: DATA = 12'b111101001111;
            14'b00_001011110001: DATA = 12'b111101010000;
            14'b00_001011110010: DATA = 12'b111101010001;
            14'b00_001011110011: DATA = 12'b111101010011;
            14'b00_001011110100: DATA = 12'b111101010100;
            14'b00_001011110101: DATA = 12'b111101010101;
            14'b00_001011110110: DATA = 12'b111101010110;
            14'b00_001011110111: DATA = 12'b111101011000;
            14'b00_001011111000: DATA = 12'b111101011001;
            14'b00_001011111001: DATA = 12'b111101011010;
            14'b00_001011111010: DATA = 12'b111101011011;
            14'b00_001011111011: DATA = 12'b111101011101;
            14'b00_001011111100: DATA = 12'b111101011110;
            14'b00_001011111101: DATA = 12'b111101011111;
            14'b00_001011111110: DATA = 12'b111101100000;
            14'b00_001011111111: DATA = 12'b111101100001;
            14'b00_001100000000: DATA = 12'b111101100011;
            14'b00_001100000001: DATA = 12'b111101100100;
            14'b00_001100000010: DATA = 12'b111101100101;
            14'b00_001100000011: DATA = 12'b111101100110;
            14'b00_001100000100: DATA = 12'b111101100111;
            14'b00_001100000101: DATA = 12'b111101101001;
            14'b00_001100000110: DATA = 12'b111101101010;
            14'b00_001100000111: DATA = 12'b111101101011;
            14'b00_001100001000: DATA = 12'b111101101100;
            14'b00_001100001001: DATA = 12'b111101101101;
            14'b00_001100001010: DATA = 12'b111101101110;
            14'b00_001100001011: DATA = 12'b111101110000;
            14'b00_001100001100: DATA = 12'b111101110001;
            14'b00_001100001101: DATA = 12'b111101110010;
            14'b00_001100001110: DATA = 12'b111101110011;
            14'b00_001100001111: DATA = 12'b111101110100;
            14'b00_001100010000: DATA = 12'b111101110101;
            14'b00_001100010001: DATA = 12'b111101110110;
            14'b00_001100010010: DATA = 12'b111101111000;
            14'b00_001100010011: DATA = 12'b111101111001;
            14'b00_001100010100: DATA = 12'b111101111010;
            14'b00_001100010101: DATA = 12'b111101111011;
            14'b00_001100010110: DATA = 12'b111101111100;
            14'b00_001100010111: DATA = 12'b111101111101;
            14'b00_001100011000: DATA = 12'b111101111110;
            14'b00_001100011001: DATA = 12'b111101111111;
            14'b00_001100011010: DATA = 12'b111110000000;
            14'b00_001100011011: DATA = 12'b111110000001;
            14'b00_001100011100: DATA = 12'b111110000011;
            14'b00_001100011101: DATA = 12'b111110000100;
            14'b00_001100011110: DATA = 12'b111110000101;
            14'b00_001100011111: DATA = 12'b111110000110;
            14'b00_001100100000: DATA = 12'b111110000111;
            14'b00_001100100001: DATA = 12'b111110001000;
            14'b00_001100100010: DATA = 12'b111110001001;
            14'b00_001100100011: DATA = 12'b111110001010;
            14'b00_001100100100: DATA = 12'b111110001011;
            14'b00_001100100101: DATA = 12'b111110001100;
            14'b00_001100100110: DATA = 12'b111110001101;
            14'b00_001100100111: DATA = 12'b111110001110;
            14'b00_001100101000: DATA = 12'b111110001111;
            14'b00_001100101001: DATA = 12'b111110010000;
            14'b00_001100101010: DATA = 12'b111110010001;
            14'b00_001100101011: DATA = 12'b111110010010;
            14'b00_001100101100: DATA = 12'b111110010011;
            14'b00_001100101101: DATA = 12'b111110010100;
            14'b00_001100101110: DATA = 12'b111110010101;
            14'b00_001100101111: DATA = 12'b111110010110;
            14'b00_001100110000: DATA = 12'b111110010111;
            14'b00_001100110001: DATA = 12'b111110011000;
            14'b00_001100110010: DATA = 12'b111110011001;
            14'b00_001100110011: DATA = 12'b111110011010;
            14'b00_001100110100: DATA = 12'b111110011011;
            14'b00_001100110101: DATA = 12'b111110011100;
            14'b00_001100110110: DATA = 12'b111110011101;
            14'b00_001100110111: DATA = 12'b111110011110;
            14'b00_001100111000: DATA = 12'b111110011111;
            14'b00_001100111001: DATA = 12'b111110100000;
            14'b00_001100111010: DATA = 12'b111110100001;
            14'b00_001100111011: DATA = 12'b111110100010;
            14'b00_001100111100: DATA = 12'b111110100011;
            14'b00_001100111101: DATA = 12'b111110100100;
            14'b00_001100111110: DATA = 12'b111110100101;
            14'b00_001100111111: DATA = 12'b111110100101;
            14'b00_001101000000: DATA = 12'b111110100110;
            14'b00_001101000001: DATA = 12'b111110100111;
            14'b00_001101000010: DATA = 12'b111110101000;
            14'b00_001101000011: DATA = 12'b111110101001;
            14'b00_001101000100: DATA = 12'b111110101010;
            14'b00_001101000101: DATA = 12'b111110101011;
            14'b00_001101000110: DATA = 12'b111110101100;
            14'b00_001101000111: DATA = 12'b111110101101;
            14'b00_001101001000: DATA = 12'b111110101110;
            14'b00_001101001001: DATA = 12'b111110101110;
            14'b00_001101001010: DATA = 12'b111110101111;
            14'b00_001101001011: DATA = 12'b111110110000;
            14'b00_001101001100: DATA = 12'b111110110001;
            14'b00_001101001101: DATA = 12'b111110110010;
            14'b00_001101001110: DATA = 12'b111110110011;
            14'b00_001101001111: DATA = 12'b111110110100;
            14'b00_001101010000: DATA = 12'b111110110100;
            14'b00_001101010001: DATA = 12'b111110110101;
            14'b00_001101010010: DATA = 12'b111110110110;
            14'b00_001101010011: DATA = 12'b111110110111;
            14'b00_001101010100: DATA = 12'b111110111000;
            14'b00_001101010101: DATA = 12'b111110111000;
            14'b00_001101010110: DATA = 12'b111110111001;
            14'b00_001101010111: DATA = 12'b111110111010;
            14'b00_001101011000: DATA = 12'b111110111011;
            14'b00_001101011001: DATA = 12'b111110111100;
            14'b00_001101011010: DATA = 12'b111110111100;
            14'b00_001101011011: DATA = 12'b111110111101;
            14'b00_001101011100: DATA = 12'b111110111110;
            14'b00_001101011101: DATA = 12'b111110111111;
            14'b00_001101011110: DATA = 12'b111111000000;
            14'b00_001101011111: DATA = 12'b111111000000;
            14'b00_001101100000: DATA = 12'b111111000001;
            14'b00_001101100001: DATA = 12'b111111000010;
            14'b00_001101100010: DATA = 12'b111111000011;
            14'b00_001101100011: DATA = 12'b111111000011;
            14'b00_001101100100: DATA = 12'b111111000100;
            14'b00_001101100101: DATA = 12'b111111000101;
            14'b00_001101100110: DATA = 12'b111111000110;
            14'b00_001101100111: DATA = 12'b111111000110;
            14'b00_001101101000: DATA = 12'b111111000111;
            14'b00_001101101001: DATA = 12'b111111001000;
            14'b00_001101101010: DATA = 12'b111111001001;
            14'b00_001101101011: DATA = 12'b111111001001;
            14'b00_001101101100: DATA = 12'b111111001010;
            14'b00_001101101101: DATA = 12'b111111001011;
            14'b00_001101101110: DATA = 12'b111111001011;
            14'b00_001101101111: DATA = 12'b111111001100;
            14'b00_001101110000: DATA = 12'b111111001101;
            14'b00_001101110001: DATA = 12'b111111001101;
            14'b00_001101110010: DATA = 12'b111111001110;
            14'b00_001101110011: DATA = 12'b111111001111;
            14'b00_001101110100: DATA = 12'b111111001111;
            14'b00_001101110101: DATA = 12'b111111010000;
            14'b00_001101110110: DATA = 12'b111111010001;
            14'b00_001101110111: DATA = 12'b111111010001;
            14'b00_001101111000: DATA = 12'b111111010010;
            14'b00_001101111001: DATA = 12'b111111010011;
            14'b00_001101111010: DATA = 12'b111111010011;
            14'b00_001101111011: DATA = 12'b111111010100;
            14'b00_001101111100: DATA = 12'b111111010101;
            14'b00_001101111101: DATA = 12'b111111010101;
            14'b00_001101111110: DATA = 12'b111111010110;
            14'b00_001101111111: DATA = 12'b111111010111;
            14'b00_001110000000: DATA = 12'b111111010111;
            14'b00_001110000001: DATA = 12'b111111011000;
            14'b00_001110000010: DATA = 12'b111111011000;
            14'b00_001110000011: DATA = 12'b111111011001;
            14'b00_001110000100: DATA = 12'b111111011010;
            14'b00_001110000101: DATA = 12'b111111011010;
            14'b00_001110000110: DATA = 12'b111111011011;
            14'b00_001110000111: DATA = 12'b111111011011;
            14'b00_001110001000: DATA = 12'b111111011100;
            14'b00_001110001001: DATA = 12'b111111011100;
            14'b00_001110001010: DATA = 12'b111111011101;
            14'b00_001110001011: DATA = 12'b111111011110;
            14'b00_001110001100: DATA = 12'b111111011110;
            14'b00_001110001101: DATA = 12'b111111011111;
            14'b00_001110001110: DATA = 12'b111111011111;
            14'b00_001110001111: DATA = 12'b111111100000;
            14'b00_001110010000: DATA = 12'b111111100000;
            14'b00_001110010001: DATA = 12'b111111100001;
            14'b00_001110010010: DATA = 12'b111111100001;
            14'b00_001110010011: DATA = 12'b111111100010;
            14'b00_001110010100: DATA = 12'b111111100010;
            14'b00_001110010101: DATA = 12'b111111100011;
            14'b00_001110010110: DATA = 12'b111111100011;
            14'b00_001110010111: DATA = 12'b111111100100;
            14'b00_001110011000: DATA = 12'b111111100101;
            14'b00_001110011001: DATA = 12'b111111100101;
            14'b00_001110011010: DATA = 12'b111111100101;
            14'b00_001110011011: DATA = 12'b111111100110;
            14'b00_001110011100: DATA = 12'b111111100110;
            14'b00_001110011101: DATA = 12'b111111100111;
            14'b00_001110011110: DATA = 12'b111111100111;
            14'b00_001110011111: DATA = 12'b111111101000;
            14'b00_001110100000: DATA = 12'b111111101000;
            14'b00_001110100001: DATA = 12'b111111101001;
            14'b00_001110100010: DATA = 12'b111111101001;
            14'b00_001110100011: DATA = 12'b111111101010;
            14'b00_001110100100: DATA = 12'b111111101010;
            14'b00_001110100101: DATA = 12'b111111101011;
            14'b00_001110100110: DATA = 12'b111111101011;
            14'b00_001110100111: DATA = 12'b111111101011;
            14'b00_001110101000: DATA = 12'b111111101100;
            14'b00_001110101001: DATA = 12'b111111101100;
            14'b00_001110101010: DATA = 12'b111111101101;
            14'b00_001110101011: DATA = 12'b111111101101;
            14'b00_001110101100: DATA = 12'b111111101110;
            14'b00_001110101101: DATA = 12'b111111101110;
            14'b00_001110101110: DATA = 12'b111111101110;
            14'b00_001110101111: DATA = 12'b111111101111;
            14'b00_001110110000: DATA = 12'b111111101111;
            14'b00_001110110001: DATA = 12'b111111101111;
            14'b00_001110110010: DATA = 12'b111111110000;
            14'b00_001110110011: DATA = 12'b111111110000;
            14'b00_001110110100: DATA = 12'b111111110001;
            14'b00_001110110101: DATA = 12'b111111110001;
            14'b00_001110110110: DATA = 12'b111111110001;
            14'b00_001110110111: DATA = 12'b111111110010;
            14'b00_001110111000: DATA = 12'b111111110010;
            14'b00_001110111001: DATA = 12'b111111110010;
            14'b00_001110111010: DATA = 12'b111111110011;
            14'b00_001110111011: DATA = 12'b111111110011;
            14'b00_001110111100: DATA = 12'b111111110011;
            14'b00_001110111101: DATA = 12'b111111110100;
            14'b00_001110111110: DATA = 12'b111111110100;
            14'b00_001110111111: DATA = 12'b111111110100;
            14'b00_001111000000: DATA = 12'b111111110101;
            14'b00_001111000001: DATA = 12'b111111110101;
            14'b00_001111000010: DATA = 12'b111111110101;
            14'b00_001111000011: DATA = 12'b111111110110;
            14'b00_001111000100: DATA = 12'b111111110110;
            14'b00_001111000101: DATA = 12'b111111110110;
            14'b00_001111000110: DATA = 12'b111111110110;
            14'b00_001111000111: DATA = 12'b111111110111;
            14'b00_001111001000: DATA = 12'b111111110111;
            14'b00_001111001001: DATA = 12'b111111110111;
            14'b00_001111001010: DATA = 12'b111111110111;
            14'b00_001111001011: DATA = 12'b111111111000;
            14'b00_001111001100: DATA = 12'b111111111000;
            14'b00_001111001101: DATA = 12'b111111111000;
            14'b00_001111001110: DATA = 12'b111111111000;
            14'b00_001111001111: DATA = 12'b111111111001;
            14'b00_001111010000: DATA = 12'b111111111001;
            14'b00_001111010001: DATA = 12'b111111111001;
            14'b00_001111010010: DATA = 12'b111111111001;
            14'b00_001111010011: DATA = 12'b111111111010;
            14'b00_001111010100: DATA = 12'b111111111010;
            14'b00_001111010101: DATA = 12'b111111111010;
            14'b00_001111010110: DATA = 12'b111111111010;
            14'b00_001111010111: DATA = 12'b111111111010;
            14'b00_001111011000: DATA = 12'b111111111011;
            14'b00_001111011001: DATA = 12'b111111111011;
            14'b00_001111011010: DATA = 12'b111111111011;
            14'b00_001111011011: DATA = 12'b111111111011;
            14'b00_001111011100: DATA = 12'b111111111011;
            14'b00_001111011101: DATA = 12'b111111111100;
            14'b00_001111011110: DATA = 12'b111111111100;
            14'b00_001111011111: DATA = 12'b111111111100;
            14'b00_001111100000: DATA = 12'b111111111100;
            14'b00_001111100001: DATA = 12'b111111111100;
            14'b00_001111100010: DATA = 12'b111111111100;
            14'b00_001111100011: DATA = 12'b111111111100;
            14'b00_001111100100: DATA = 12'b111111111101;
            14'b00_001111100101: DATA = 12'b111111111101;
            14'b00_001111100110: DATA = 12'b111111111101;
            14'b00_001111100111: DATA = 12'b111111111101;
            14'b00_001111101000: DATA = 12'b111111111101;
            14'b00_001111101001: DATA = 12'b111111111101;
            14'b00_001111101010: DATA = 12'b111111111101;
            14'b00_001111101011: DATA = 12'b111111111101;
            14'b00_001111101100: DATA = 12'b111111111110;
            14'b00_001111101101: DATA = 12'b111111111110;
            14'b00_001111101110: DATA = 12'b111111111110;
            14'b00_001111101111: DATA = 12'b111111111110;
            14'b00_001111110000: DATA = 12'b111111111110;
            14'b00_001111110001: DATA = 12'b111111111110;
            14'b00_001111110010: DATA = 12'b111111111110;
            14'b00_001111110011: DATA = 12'b111111111110;
            14'b00_001111110100: DATA = 12'b111111111110;
            14'b00_001111110101: DATA = 12'b111111111110;
            14'b00_001111110110: DATA = 12'b111111111110;
            14'b00_001111110111: DATA = 12'b111111111110;
            14'b00_001111111000: DATA = 12'b111111111110;
            14'b00_001111111001: DATA = 12'b111111111110;
            14'b00_001111111010: DATA = 12'b111111111110;
            14'b00_001111111011: DATA = 12'b111111111110;
            14'b00_001111111100: DATA = 12'b111111111110;
            14'b00_001111111101: DATA = 12'b111111111110;
            14'b00_001111111110: DATA = 12'b111111111110;
            14'b00_001111111111: DATA = 12'b111111111110;
            14'b00_010000000000: DATA = 12'b111111111111;
            14'b00_010000000001: DATA = 12'b111111111110;
            14'b00_010000000010: DATA = 12'b111111111110;
            14'b00_010000000011: DATA = 12'b111111111110;
            14'b00_010000000100: DATA = 12'b111111111110;
            14'b00_010000000101: DATA = 12'b111111111110;
            14'b00_010000000110: DATA = 12'b111111111110;
            14'b00_010000000111: DATA = 12'b111111111110;
            14'b00_010000001000: DATA = 12'b111111111110;
            14'b00_010000001001: DATA = 12'b111111111110;
            14'b00_010000001010: DATA = 12'b111111111110;
            14'b00_010000001011: DATA = 12'b111111111110;
            14'b00_010000001100: DATA = 12'b111111111110;
            14'b00_010000001101: DATA = 12'b111111111110;
            14'b00_010000001110: DATA = 12'b111111111110;
            14'b00_010000001111: DATA = 12'b111111111110;
            14'b00_010000010000: DATA = 12'b111111111110;
            14'b00_010000010001: DATA = 12'b111111111110;
            14'b00_010000010010: DATA = 12'b111111111110;
            14'b00_010000010011: DATA = 12'b111111111110;
            14'b00_010000010100: DATA = 12'b111111111110;
            14'b00_010000010101: DATA = 12'b111111111101;
            14'b00_010000010110: DATA = 12'b111111111101;
            14'b00_010000010111: DATA = 12'b111111111101;
            14'b00_010000011000: DATA = 12'b111111111101;
            14'b00_010000011001: DATA = 12'b111111111101;
            14'b00_010000011010: DATA = 12'b111111111101;
            14'b00_010000011011: DATA = 12'b111111111101;
            14'b00_010000011100: DATA = 12'b111111111101;
            14'b00_010000011101: DATA = 12'b111111111100;
            14'b00_010000011110: DATA = 12'b111111111100;
            14'b00_010000011111: DATA = 12'b111111111100;
            14'b00_010000100000: DATA = 12'b111111111100;
            14'b00_010000100001: DATA = 12'b111111111100;
            14'b00_010000100010: DATA = 12'b111111111100;
            14'b00_010000100011: DATA = 12'b111111111100;
            14'b00_010000100100: DATA = 12'b111111111011;
            14'b00_010000100101: DATA = 12'b111111111011;
            14'b00_010000100110: DATA = 12'b111111111011;
            14'b00_010000100111: DATA = 12'b111111111011;
            14'b00_010000101000: DATA = 12'b111111111011;
            14'b00_010000101001: DATA = 12'b111111111010;
            14'b00_010000101010: DATA = 12'b111111111010;
            14'b00_010000101011: DATA = 12'b111111111010;
            14'b00_010000101100: DATA = 12'b111111111010;
            14'b00_010000101101: DATA = 12'b111111111010;
            14'b00_010000101110: DATA = 12'b111111111001;
            14'b00_010000101111: DATA = 12'b111111111001;
            14'b00_010000110000: DATA = 12'b111111111001;
            14'b00_010000110001: DATA = 12'b111111111001;
            14'b00_010000110010: DATA = 12'b111111111000;
            14'b00_010000110011: DATA = 12'b111111111000;
            14'b00_010000110100: DATA = 12'b111111111000;
            14'b00_010000110101: DATA = 12'b111111111000;
            14'b00_010000110110: DATA = 12'b111111110111;
            14'b00_010000110111: DATA = 12'b111111110111;
            14'b00_010000111000: DATA = 12'b111111110111;
            14'b00_010000111001: DATA = 12'b111111110111;
            14'b00_010000111010: DATA = 12'b111111110110;
            14'b00_010000111011: DATA = 12'b111111110110;
            14'b00_010000111100: DATA = 12'b111111110110;
            14'b00_010000111101: DATA = 12'b111111110110;
            14'b00_010000111110: DATA = 12'b111111110101;
            14'b00_010000111111: DATA = 12'b111111110101;
            14'b00_010001000000: DATA = 12'b111111110101;
            14'b00_010001000001: DATA = 12'b111111110100;
            14'b00_010001000010: DATA = 12'b111111110100;
            14'b00_010001000011: DATA = 12'b111111110100;
            14'b00_010001000100: DATA = 12'b111111110011;
            14'b00_010001000101: DATA = 12'b111111110011;
            14'b00_010001000110: DATA = 12'b111111110011;
            14'b00_010001000111: DATA = 12'b111111110010;
            14'b00_010001001000: DATA = 12'b111111110010;
            14'b00_010001001001: DATA = 12'b111111110010;
            14'b00_010001001010: DATA = 12'b111111110001;
            14'b00_010001001011: DATA = 12'b111111110001;
            14'b00_010001001100: DATA = 12'b111111110001;
            14'b00_010001001101: DATA = 12'b111111110000;
            14'b00_010001001110: DATA = 12'b111111110000;
            14'b00_010001001111: DATA = 12'b111111101111;
            14'b00_010001010000: DATA = 12'b111111101111;
            14'b00_010001010001: DATA = 12'b111111101111;
            14'b00_010001010010: DATA = 12'b111111101110;
            14'b00_010001010011: DATA = 12'b111111101110;
            14'b00_010001010100: DATA = 12'b111111101110;
            14'b00_010001010101: DATA = 12'b111111101101;
            14'b00_010001010110: DATA = 12'b111111101101;
            14'b00_010001010111: DATA = 12'b111111101100;
            14'b00_010001011000: DATA = 12'b111111101100;
            14'b00_010001011001: DATA = 12'b111111101011;
            14'b00_010001011010: DATA = 12'b111111101011;
            14'b00_010001011011: DATA = 12'b111111101011;
            14'b00_010001011100: DATA = 12'b111111101010;
            14'b00_010001011101: DATA = 12'b111111101010;
            14'b00_010001011110: DATA = 12'b111111101001;
            14'b00_010001011111: DATA = 12'b111111101001;
            14'b00_010001100000: DATA = 12'b111111101000;
            14'b00_010001100001: DATA = 12'b111111101000;
            14'b00_010001100010: DATA = 12'b111111100111;
            14'b00_010001100011: DATA = 12'b111111100111;
            14'b00_010001100100: DATA = 12'b111111100110;
            14'b00_010001100101: DATA = 12'b111111100110;
            14'b00_010001100110: DATA = 12'b111111100101;
            14'b00_010001100111: DATA = 12'b111111100101;
            14'b00_010001101000: DATA = 12'b111111100101;
            14'b00_010001101001: DATA = 12'b111111100100;
            14'b00_010001101010: DATA = 12'b111111100011;
            14'b00_010001101011: DATA = 12'b111111100011;
            14'b00_010001101100: DATA = 12'b111111100010;
            14'b00_010001101101: DATA = 12'b111111100010;
            14'b00_010001101110: DATA = 12'b111111100001;
            14'b00_010001101111: DATA = 12'b111111100001;
            14'b00_010001110000: DATA = 12'b111111100000;
            14'b00_010001110001: DATA = 12'b111111100000;
            14'b00_010001110010: DATA = 12'b111111011111;
            14'b00_010001110011: DATA = 12'b111111011111;
            14'b00_010001110100: DATA = 12'b111111011110;
            14'b00_010001110101: DATA = 12'b111111011110;
            14'b00_010001110110: DATA = 12'b111111011101;
            14'b00_010001110111: DATA = 12'b111111011100;
            14'b00_010001111000: DATA = 12'b111111011100;
            14'b00_010001111001: DATA = 12'b111111011011;
            14'b00_010001111010: DATA = 12'b111111011011;
            14'b00_010001111011: DATA = 12'b111111011010;
            14'b00_010001111100: DATA = 12'b111111011010;
            14'b00_010001111101: DATA = 12'b111111011001;
            14'b00_010001111110: DATA = 12'b111111011000;
            14'b00_010001111111: DATA = 12'b111111011000;
            14'b00_010010000000: DATA = 12'b111111010111;
            14'b00_010010000001: DATA = 12'b111111010111;
            14'b00_010010000010: DATA = 12'b111111010110;
            14'b00_010010000011: DATA = 12'b111111010101;
            14'b00_010010000100: DATA = 12'b111111010101;
            14'b00_010010000101: DATA = 12'b111111010100;
            14'b00_010010000110: DATA = 12'b111111010011;
            14'b00_010010000111: DATA = 12'b111111010011;
            14'b00_010010001000: DATA = 12'b111111010010;
            14'b00_010010001001: DATA = 12'b111111010001;
            14'b00_010010001010: DATA = 12'b111111010001;
            14'b00_010010001011: DATA = 12'b111111010000;
            14'b00_010010001100: DATA = 12'b111111001111;
            14'b00_010010001101: DATA = 12'b111111001111;
            14'b00_010010001110: DATA = 12'b111111001110;
            14'b00_010010001111: DATA = 12'b111111001101;
            14'b00_010010010000: DATA = 12'b111111001101;
            14'b00_010010010001: DATA = 12'b111111001100;
            14'b00_010010010010: DATA = 12'b111111001011;
            14'b00_010010010011: DATA = 12'b111111001011;
            14'b00_010010010100: DATA = 12'b111111001010;
            14'b00_010010010101: DATA = 12'b111111001001;
            14'b00_010010010110: DATA = 12'b111111001001;
            14'b00_010010010111: DATA = 12'b111111001000;
            14'b00_010010011000: DATA = 12'b111111000111;
            14'b00_010010011001: DATA = 12'b111111000110;
            14'b00_010010011010: DATA = 12'b111111000110;
            14'b00_010010011011: DATA = 12'b111111000101;
            14'b00_010010011100: DATA = 12'b111111000100;
            14'b00_010010011101: DATA = 12'b111111000011;
            14'b00_010010011110: DATA = 12'b111111000011;
            14'b00_010010011111: DATA = 12'b111111000010;
            14'b00_010010100000: DATA = 12'b111111000001;
            14'b00_010010100001: DATA = 12'b111111000000;
            14'b00_010010100010: DATA = 12'b111111000000;
            14'b00_010010100011: DATA = 12'b111110111111;
            14'b00_010010100100: DATA = 12'b111110111110;
            14'b00_010010100101: DATA = 12'b111110111101;
            14'b00_010010100110: DATA = 12'b111110111100;
            14'b00_010010100111: DATA = 12'b111110111100;
            14'b00_010010101000: DATA = 12'b111110111011;
            14'b00_010010101001: DATA = 12'b111110111010;
            14'b00_010010101010: DATA = 12'b111110111001;
            14'b00_010010101011: DATA = 12'b111110111000;
            14'b00_010010101100: DATA = 12'b111110111000;
            14'b00_010010101101: DATA = 12'b111110110111;
            14'b00_010010101110: DATA = 12'b111110110110;
            14'b00_010010101111: DATA = 12'b111110110101;
            14'b00_010010110000: DATA = 12'b111110110100;
            14'b00_010010110001: DATA = 12'b111110110100;
            14'b00_010010110010: DATA = 12'b111110110011;
            14'b00_010010110011: DATA = 12'b111110110010;
            14'b00_010010110100: DATA = 12'b111110110001;
            14'b00_010010110101: DATA = 12'b111110110000;
            14'b00_010010110110: DATA = 12'b111110101111;
            14'b00_010010110111: DATA = 12'b111110101110;
            14'b00_010010111000: DATA = 12'b111110101110;
            14'b00_010010111001: DATA = 12'b111110101101;
            14'b00_010010111010: DATA = 12'b111110101100;
            14'b00_010010111011: DATA = 12'b111110101011;
            14'b00_010010111100: DATA = 12'b111110101010;
            14'b00_010010111101: DATA = 12'b111110101001;
            14'b00_010010111110: DATA = 12'b111110101000;
            14'b00_010010111111: DATA = 12'b111110100111;
            14'b00_010011000000: DATA = 12'b111110100110;
            14'b00_010011000001: DATA = 12'b111110100101;
            14'b00_010011000010: DATA = 12'b111110100101;
            14'b00_010011000011: DATA = 12'b111110100100;
            14'b00_010011000100: DATA = 12'b111110100011;
            14'b00_010011000101: DATA = 12'b111110100010;
            14'b00_010011000110: DATA = 12'b111110100001;
            14'b00_010011000111: DATA = 12'b111110100000;
            14'b00_010011001000: DATA = 12'b111110011111;
            14'b00_010011001001: DATA = 12'b111110011110;
            14'b00_010011001010: DATA = 12'b111110011101;
            14'b00_010011001011: DATA = 12'b111110011100;
            14'b00_010011001100: DATA = 12'b111110011011;
            14'b00_010011001101: DATA = 12'b111110011010;
            14'b00_010011001110: DATA = 12'b111110011001;
            14'b00_010011001111: DATA = 12'b111110011000;
            14'b00_010011010000: DATA = 12'b111110010111;
            14'b00_010011010001: DATA = 12'b111110010110;
            14'b00_010011010010: DATA = 12'b111110010101;
            14'b00_010011010011: DATA = 12'b111110010100;
            14'b00_010011010100: DATA = 12'b111110010011;
            14'b00_010011010101: DATA = 12'b111110010010;
            14'b00_010011010110: DATA = 12'b111110010001;
            14'b00_010011010111: DATA = 12'b111110010000;
            14'b00_010011011000: DATA = 12'b111110001111;
            14'b00_010011011001: DATA = 12'b111110001110;
            14'b00_010011011010: DATA = 12'b111110001101;
            14'b00_010011011011: DATA = 12'b111110001100;
            14'b00_010011011100: DATA = 12'b111110001011;
            14'b00_010011011101: DATA = 12'b111110001010;
            14'b00_010011011110: DATA = 12'b111110001001;
            14'b00_010011011111: DATA = 12'b111110001000;
            14'b00_010011100000: DATA = 12'b111110000111;
            14'b00_010011100001: DATA = 12'b111110000110;
            14'b00_010011100010: DATA = 12'b111110000101;
            14'b00_010011100011: DATA = 12'b111110000100;
            14'b00_010011100100: DATA = 12'b111110000011;
            14'b00_010011100101: DATA = 12'b111110000001;
            14'b00_010011100110: DATA = 12'b111110000000;
            14'b00_010011100111: DATA = 12'b111101111111;
            14'b00_010011101000: DATA = 12'b111101111110;
            14'b00_010011101001: DATA = 12'b111101111101;
            14'b00_010011101010: DATA = 12'b111101111100;
            14'b00_010011101011: DATA = 12'b111101111011;
            14'b00_010011101100: DATA = 12'b111101111010;
            14'b00_010011101101: DATA = 12'b111101111001;
            14'b00_010011101110: DATA = 12'b111101111000;
            14'b00_010011101111: DATA = 12'b111101110110;
            14'b00_010011110000: DATA = 12'b111101110101;
            14'b00_010011110001: DATA = 12'b111101110100;
            14'b00_010011110010: DATA = 12'b111101110011;
            14'b00_010011110011: DATA = 12'b111101110010;
            14'b00_010011110100: DATA = 12'b111101110001;
            14'b00_010011110101: DATA = 12'b111101110000;
            14'b00_010011110110: DATA = 12'b111101101110;
            14'b00_010011110111: DATA = 12'b111101101101;
            14'b00_010011111000: DATA = 12'b111101101100;
            14'b00_010011111001: DATA = 12'b111101101011;
            14'b00_010011111010: DATA = 12'b111101101010;
            14'b00_010011111011: DATA = 12'b111101101001;
            14'b00_010011111100: DATA = 12'b111101100111;
            14'b00_010011111101: DATA = 12'b111101100110;
            14'b00_010011111110: DATA = 12'b111101100101;
            14'b00_010011111111: DATA = 12'b111101100100;
            14'b00_010100000000: DATA = 12'b111101100011;
            14'b00_010100000001: DATA = 12'b111101100001;
            14'b00_010100000010: DATA = 12'b111101100000;
            14'b00_010100000011: DATA = 12'b111101011111;
            14'b00_010100000100: DATA = 12'b111101011110;
            14'b00_010100000101: DATA = 12'b111101011101;
            14'b00_010100000110: DATA = 12'b111101011011;
            14'b00_010100000111: DATA = 12'b111101011010;
            14'b00_010100001000: DATA = 12'b111101011001;
            14'b00_010100001001: DATA = 12'b111101011000;
            14'b00_010100001010: DATA = 12'b111101010110;
            14'b00_010100001011: DATA = 12'b111101010101;
            14'b00_010100001100: DATA = 12'b111101010100;
            14'b00_010100001101: DATA = 12'b111101010011;
            14'b00_010100001110: DATA = 12'b111101010001;
            14'b00_010100001111: DATA = 12'b111101010000;
            14'b00_010100010000: DATA = 12'b111101001111;
            14'b00_010100010001: DATA = 12'b111101001110;
            14'b00_010100010010: DATA = 12'b111101001100;
            14'b00_010100010011: DATA = 12'b111101001011;
            14'b00_010100010100: DATA = 12'b111101001010;
            14'b00_010100010101: DATA = 12'b111101001000;
            14'b00_010100010110: DATA = 12'b111101000111;
            14'b00_010100010111: DATA = 12'b111101000110;
            14'b00_010100011000: DATA = 12'b111101000101;
            14'b00_010100011001: DATA = 12'b111101000011;
            14'b00_010100011010: DATA = 12'b111101000010;
            14'b00_010100011011: DATA = 12'b111101000001;
            14'b00_010100011100: DATA = 12'b111100111111;
            14'b00_010100011101: DATA = 12'b111100111110;
            14'b00_010100011110: DATA = 12'b111100111101;
            14'b00_010100011111: DATA = 12'b111100111011;
            14'b00_010100100000: DATA = 12'b111100111010;
            14'b00_010100100001: DATA = 12'b111100111001;
            14'b00_010100100010: DATA = 12'b111100110111;
            14'b00_010100100011: DATA = 12'b111100110110;
            14'b00_010100100100: DATA = 12'b111100110101;
            14'b00_010100100101: DATA = 12'b111100110011;
            14'b00_010100100110: DATA = 12'b111100110010;
            14'b00_010100100111: DATA = 12'b111100110000;
            14'b00_010100101000: DATA = 12'b111100101111;
            14'b00_010100101001: DATA = 12'b111100101110;
            14'b00_010100101010: DATA = 12'b111100101100;
            14'b00_010100101011: DATA = 12'b111100101011;
            14'b00_010100101100: DATA = 12'b111100101010;
            14'b00_010100101101: DATA = 12'b111100101000;
            14'b00_010100101110: DATA = 12'b111100100111;
            14'b00_010100101111: DATA = 12'b111100100101;
            14'b00_010100110000: DATA = 12'b111100100100;
            14'b00_010100110001: DATA = 12'b111100100011;
            14'b00_010100110010: DATA = 12'b111100100001;
            14'b00_010100110011: DATA = 12'b111100100000;
            14'b00_010100110100: DATA = 12'b111100011110;
            14'b00_010100110101: DATA = 12'b111100011101;
            14'b00_010100110110: DATA = 12'b111100011011;
            14'b00_010100110111: DATA = 12'b111100011010;
            14'b00_010100111000: DATA = 12'b111100011000;
            14'b00_010100111001: DATA = 12'b111100010111;
            14'b00_010100111010: DATA = 12'b111100010110;
            14'b00_010100111011: DATA = 12'b111100010100;
            14'b00_010100111100: DATA = 12'b111100010011;
            14'b00_010100111101: DATA = 12'b111100010001;
            14'b00_010100111110: DATA = 12'b111100010000;
            14'b00_010100111111: DATA = 12'b111100001110;
            14'b00_010101000000: DATA = 12'b111100001101;
            14'b00_010101000001: DATA = 12'b111100001011;
            14'b00_010101000010: DATA = 12'b111100001010;
            14'b00_010101000011: DATA = 12'b111100001000;
            14'b00_010101000100: DATA = 12'b111100000111;
            14'b00_010101000101: DATA = 12'b111100000101;
            14'b00_010101000110: DATA = 12'b111100000100;
            14'b00_010101000111: DATA = 12'b111100000010;
            14'b00_010101001000: DATA = 12'b111100000001;
            14'b00_010101001001: DATA = 12'b111011111111;
            14'b00_010101001010: DATA = 12'b111011111110;
            14'b00_010101001011: DATA = 12'b111011111100;
            14'b00_010101001100: DATA = 12'b111011111011;
            14'b00_010101001101: DATA = 12'b111011111001;
            14'b00_010101001110: DATA = 12'b111011111000;
            14'b00_010101001111: DATA = 12'b111011110110;
            14'b00_010101010000: DATA = 12'b111011110101;
            14'b00_010101010001: DATA = 12'b111011110011;
            14'b00_010101010010: DATA = 12'b111011110001;
            14'b00_010101010011: DATA = 12'b111011110000;
            14'b00_010101010100: DATA = 12'b111011101110;
            14'b00_010101010101: DATA = 12'b111011101101;
            14'b00_010101010110: DATA = 12'b111011101011;
            14'b00_010101010111: DATA = 12'b111011101010;
            14'b00_010101011000: DATA = 12'b111011101000;
            14'b00_010101011001: DATA = 12'b111011100110;
            14'b00_010101011010: DATA = 12'b111011100101;
            14'b00_010101011011: DATA = 12'b111011100011;
            14'b00_010101011100: DATA = 12'b111011100010;
            14'b00_010101011101: DATA = 12'b111011100000;
            14'b00_010101011110: DATA = 12'b111011011110;
            14'b00_010101011111: DATA = 12'b111011011101;
            14'b00_010101100000: DATA = 12'b111011011011;
            14'b00_010101100001: DATA = 12'b111011011010;
            14'b00_010101100010: DATA = 12'b111011011000;
            14'b00_010101100011: DATA = 12'b111011010110;
            14'b00_010101100100: DATA = 12'b111011010101;
            14'b00_010101100101: DATA = 12'b111011010011;
            14'b00_010101100110: DATA = 12'b111011010010;
            14'b00_010101100111: DATA = 12'b111011010000;
            14'b00_010101101000: DATA = 12'b111011001110;
            14'b00_010101101001: DATA = 12'b111011001101;
            14'b00_010101101010: DATA = 12'b111011001011;
            14'b00_010101101011: DATA = 12'b111011001001;
            14'b00_010101101100: DATA = 12'b111011001000;
            14'b00_010101101101: DATA = 12'b111011000110;
            14'b00_010101101110: DATA = 12'b111011000100;
            14'b00_010101101111: DATA = 12'b111011000011;
            14'b00_010101110000: DATA = 12'b111011000001;
            14'b00_010101110001: DATA = 12'b111010111111;
            14'b00_010101110010: DATA = 12'b111010111110;
            14'b00_010101110011: DATA = 12'b111010111100;
            14'b00_010101110100: DATA = 12'b111010111010;
            14'b00_010101110101: DATA = 12'b111010111000;
            14'b00_010101110110: DATA = 12'b111010110111;
            14'b00_010101110111: DATA = 12'b111010110101;
            14'b00_010101111000: DATA = 12'b111010110011;
            14'b00_010101111001: DATA = 12'b111010110010;
            14'b00_010101111010: DATA = 12'b111010110000;
            14'b00_010101111011: DATA = 12'b111010101110;
            14'b00_010101111100: DATA = 12'b111010101100;
            14'b00_010101111101: DATA = 12'b111010101011;
            14'b00_010101111110: DATA = 12'b111010101001;
            14'b00_010101111111: DATA = 12'b111010100111;
            14'b00_010110000000: DATA = 12'b111010100110;
            14'b00_010110000001: DATA = 12'b111010100100;
            14'b00_010110000010: DATA = 12'b111010100010;
            14'b00_010110000011: DATA = 12'b111010100000;
            14'b00_010110000100: DATA = 12'b111010011111;
            14'b00_010110000101: DATA = 12'b111010011101;
            14'b00_010110000110: DATA = 12'b111010011011;
            14'b00_010110000111: DATA = 12'b111010011001;
            14'b00_010110001000: DATA = 12'b111010010111;
            14'b00_010110001001: DATA = 12'b111010010110;
            14'b00_010110001010: DATA = 12'b111010010100;
            14'b00_010110001011: DATA = 12'b111010010010;
            14'b00_010110001100: DATA = 12'b111010010000;
            14'b00_010110001101: DATA = 12'b111010001111;
            14'b00_010110001110: DATA = 12'b111010001101;
            14'b00_010110001111: DATA = 12'b111010001011;
            14'b00_010110010000: DATA = 12'b111010001001;
            14'b00_010110010001: DATA = 12'b111010000111;
            14'b00_010110010010: DATA = 12'b111010000101;
            14'b00_010110010011: DATA = 12'b111010000100;
            14'b00_010110010100: DATA = 12'b111010000010;
            14'b00_010110010101: DATA = 12'b111010000000;
            14'b00_010110010110: DATA = 12'b111001111110;
            14'b00_010110010111: DATA = 12'b111001111100;
            14'b00_010110011000: DATA = 12'b111001111011;
            14'b00_010110011001: DATA = 12'b111001111001;
            14'b00_010110011010: DATA = 12'b111001110111;
            14'b00_010110011011: DATA = 12'b111001110101;
            14'b00_010110011100: DATA = 12'b111001110011;
            14'b00_010110011101: DATA = 12'b111001110001;
            14'b00_010110011110: DATA = 12'b111001101111;
            14'b00_010110011111: DATA = 12'b111001101110;
            14'b00_010110100000: DATA = 12'b111001101100;
            14'b00_010110100001: DATA = 12'b111001101010;
            14'b00_010110100010: DATA = 12'b111001101000;
            14'b00_010110100011: DATA = 12'b111001100110;
            14'b00_010110100100: DATA = 12'b111001100100;
            14'b00_010110100101: DATA = 12'b111001100010;
            14'b00_010110100110: DATA = 12'b111001100000;
            14'b00_010110100111: DATA = 12'b111001011110;
            14'b00_010110101000: DATA = 12'b111001011101;
            14'b00_010110101001: DATA = 12'b111001011011;
            14'b00_010110101010: DATA = 12'b111001011001;
            14'b00_010110101011: DATA = 12'b111001010111;
            14'b00_010110101100: DATA = 12'b111001010101;
            14'b00_010110101101: DATA = 12'b111001010011;
            14'b00_010110101110: DATA = 12'b111001010001;
            14'b00_010110101111: DATA = 12'b111001001111;
            14'b00_010110110000: DATA = 12'b111001001101;
            14'b00_010110110001: DATA = 12'b111001001011;
            14'b00_010110110010: DATA = 12'b111001001001;
            14'b00_010110110011: DATA = 12'b111001000111;
            14'b00_010110110100: DATA = 12'b111001000101;
            14'b00_010110110101: DATA = 12'b111001000100;
            14'b00_010110110110: DATA = 12'b111001000010;
            14'b00_010110110111: DATA = 12'b111001000000;
            14'b00_010110111000: DATA = 12'b111000111110;
            14'b00_010110111001: DATA = 12'b111000111100;
            14'b00_010110111010: DATA = 12'b111000111010;
            14'b00_010110111011: DATA = 12'b111000111000;
            14'b00_010110111100: DATA = 12'b111000110110;
            14'b00_010110111101: DATA = 12'b111000110100;
            14'b00_010110111110: DATA = 12'b111000110010;
            14'b00_010110111111: DATA = 12'b111000110000;
            14'b00_010111000000: DATA = 12'b111000101110;
            14'b00_010111000001: DATA = 12'b111000101100;
            14'b00_010111000010: DATA = 12'b111000101010;
            14'b00_010111000011: DATA = 12'b111000101000;
            14'b00_010111000100: DATA = 12'b111000100110;
            14'b00_010111000101: DATA = 12'b111000100100;
            14'b00_010111000110: DATA = 12'b111000100010;
            14'b00_010111000111: DATA = 12'b111000100000;
            14'b00_010111001000: DATA = 12'b111000011110;
            14'b00_010111001001: DATA = 12'b111000011100;
            14'b00_010111001010: DATA = 12'b111000011010;
            14'b00_010111001011: DATA = 12'b111000011000;
            14'b00_010111001100: DATA = 12'b111000010110;
            14'b00_010111001101: DATA = 12'b111000010100;
            14'b00_010111001110: DATA = 12'b111000010010;
            14'b00_010111001111: DATA = 12'b111000010000;
            14'b00_010111010000: DATA = 12'b111000001110;
            14'b00_010111010001: DATA = 12'b111000001011;
            14'b00_010111010010: DATA = 12'b111000001001;
            14'b00_010111010011: DATA = 12'b111000000111;
            14'b00_010111010100: DATA = 12'b111000000101;
            14'b00_010111010101: DATA = 12'b111000000011;
            14'b00_010111010110: DATA = 12'b111000000001;
            14'b00_010111010111: DATA = 12'b110111111111;
            14'b00_010111011000: DATA = 12'b110111111101;
            14'b00_010111011001: DATA = 12'b110111111011;
            14'b00_010111011010: DATA = 12'b110111111001;
            14'b00_010111011011: DATA = 12'b110111110111;
            14'b00_010111011100: DATA = 12'b110111110101;
            14'b00_010111011101: DATA = 12'b110111110011;
            14'b00_010111011110: DATA = 12'b110111110000;
            14'b00_010111011111: DATA = 12'b110111101110;
            14'b00_010111100000: DATA = 12'b110111101100;
            14'b00_010111100001: DATA = 12'b110111101010;
            14'b00_010111100010: DATA = 12'b110111101000;
            14'b00_010111100011: DATA = 12'b110111100110;
            14'b00_010111100100: DATA = 12'b110111100100;
            14'b00_010111100101: DATA = 12'b110111100010;
            14'b00_010111100110: DATA = 12'b110111100000;
            14'b00_010111100111: DATA = 12'b110111011101;
            14'b00_010111101000: DATA = 12'b110111011011;
            14'b00_010111101001: DATA = 12'b110111011001;
            14'b00_010111101010: DATA = 12'b110111010111;
            14'b00_010111101011: DATA = 12'b110111010101;
            14'b00_010111101100: DATA = 12'b110111010011;
            14'b00_010111101101: DATA = 12'b110111010001;
            14'b00_010111101110: DATA = 12'b110111001110;
            14'b00_010111101111: DATA = 12'b110111001100;
            14'b00_010111110000: DATA = 12'b110111001010;
            14'b00_010111110001: DATA = 12'b110111001000;
            14'b00_010111110010: DATA = 12'b110111000110;
            14'b00_010111110011: DATA = 12'b110111000100;
            14'b00_010111110100: DATA = 12'b110111000001;
            14'b00_010111110101: DATA = 12'b110110111111;
            14'b00_010111110110: DATA = 12'b110110111101;
            14'b00_010111110111: DATA = 12'b110110111011;
            14'b00_010111111000: DATA = 12'b110110111001;
            14'b00_010111111001: DATA = 12'b110110110110;
            14'b00_010111111010: DATA = 12'b110110110100;
            14'b00_010111111011: DATA = 12'b110110110010;
            14'b00_010111111100: DATA = 12'b110110110000;
            14'b00_010111111101: DATA = 12'b110110101110;
            14'b00_010111111110: DATA = 12'b110110101011;
            14'b00_010111111111: DATA = 12'b110110101001;
            14'b00_011000000000: DATA = 12'b110110100111;
            14'b00_011000000001: DATA = 12'b110110100101;
            14'b00_011000000010: DATA = 12'b110110100011;
            14'b00_011000000011: DATA = 12'b110110100000;
            14'b00_011000000100: DATA = 12'b110110011110;
            14'b00_011000000101: DATA = 12'b110110011100;
            14'b00_011000000110: DATA = 12'b110110011010;
            14'b00_011000000111: DATA = 12'b110110010111;
            14'b00_011000001000: DATA = 12'b110110010101;
            14'b00_011000001001: DATA = 12'b110110010011;
            14'b00_011000001010: DATA = 12'b110110010001;
            14'b00_011000001011: DATA = 12'b110110001110;
            14'b00_011000001100: DATA = 12'b110110001100;
            14'b00_011000001101: DATA = 12'b110110001010;
            14'b00_011000001110: DATA = 12'b110110001000;
            14'b00_011000001111: DATA = 12'b110110000101;
            14'b00_011000010000: DATA = 12'b110110000011;
            14'b00_011000010001: DATA = 12'b110110000001;
            14'b00_011000010010: DATA = 12'b110101111110;
            14'b00_011000010011: DATA = 12'b110101111100;
            14'b00_011000010100: DATA = 12'b110101111010;
            14'b00_011000010101: DATA = 12'b110101111000;
            14'b00_011000010110: DATA = 12'b110101110101;
            14'b00_011000010111: DATA = 12'b110101110011;
            14'b00_011000011000: DATA = 12'b110101110001;
            14'b00_011000011001: DATA = 12'b110101101110;
            14'b00_011000011010: DATA = 12'b110101101100;
            14'b00_011000011011: DATA = 12'b110101101010;
            14'b00_011000011100: DATA = 12'b110101100111;
            14'b00_011000011101: DATA = 12'b110101100101;
            14'b00_011000011110: DATA = 12'b110101100011;
            14'b00_011000011111: DATA = 12'b110101100001;
            14'b00_011000100000: DATA = 12'b110101011110;
            14'b00_011000100001: DATA = 12'b110101011100;
            14'b00_011000100010: DATA = 12'b110101011010;
            14'b00_011000100011: DATA = 12'b110101010111;
            14'b00_011000100100: DATA = 12'b110101010101;
            14'b00_011000100101: DATA = 12'b110101010011;
            14'b00_011000100110: DATA = 12'b110101010000;
            14'b00_011000100111: DATA = 12'b110101001110;
            14'b00_011000101000: DATA = 12'b110101001011;
            14'b00_011000101001: DATA = 12'b110101001001;
            14'b00_011000101010: DATA = 12'b110101000111;
            14'b00_011000101011: DATA = 12'b110101000100;
            14'b00_011000101100: DATA = 12'b110101000010;
            14'b00_011000101101: DATA = 12'b110101000000;
            14'b00_011000101110: DATA = 12'b110100111101;
            14'b00_011000101111: DATA = 12'b110100111011;
            14'b00_011000110000: DATA = 12'b110100111001;
            14'b00_011000110001: DATA = 12'b110100110110;
            14'b00_011000110010: DATA = 12'b110100110100;
            14'b00_011000110011: DATA = 12'b110100110001;
            14'b00_011000110100: DATA = 12'b110100101111;
            14'b00_011000110101: DATA = 12'b110100101101;
            14'b00_011000110110: DATA = 12'b110100101010;
            14'b00_011000110111: DATA = 12'b110100101000;
            14'b00_011000111000: DATA = 12'b110100100101;
            14'b00_011000111001: DATA = 12'b110100100011;
            14'b00_011000111010: DATA = 12'b110100100001;
            14'b00_011000111011: DATA = 12'b110100011110;
            14'b00_011000111100: DATA = 12'b110100011100;
            14'b00_011000111101: DATA = 12'b110100011001;
            14'b00_011000111110: DATA = 12'b110100010111;
            14'b00_011000111111: DATA = 12'b110100010101;
            14'b00_011001000000: DATA = 12'b110100010010;
            14'b00_011001000001: DATA = 12'b110100010000;
            14'b00_011001000010: DATA = 12'b110100001101;
            14'b00_011001000011: DATA = 12'b110100001011;
            14'b00_011001000100: DATA = 12'b110100001000;
            14'b00_011001000101: DATA = 12'b110100000110;
            14'b00_011001000110: DATA = 12'b110100000011;
            14'b00_011001000111: DATA = 12'b110100000001;
            14'b00_011001001000: DATA = 12'b110011111111;
            14'b00_011001001001: DATA = 12'b110011111100;
            14'b00_011001001010: DATA = 12'b110011111010;
            14'b00_011001001011: DATA = 12'b110011110111;
            14'b00_011001001100: DATA = 12'b110011110101;
            14'b00_011001001101: DATA = 12'b110011110010;
            14'b00_011001001110: DATA = 12'b110011110000;
            14'b00_011001001111: DATA = 12'b110011101101;
            14'b00_011001010000: DATA = 12'b110011101011;
            14'b00_011001010001: DATA = 12'b110011101000;
            14'b00_011001010010: DATA = 12'b110011100110;
            14'b00_011001010011: DATA = 12'b110011100011;
            14'b00_011001010100: DATA = 12'b110011100001;
            14'b00_011001010101: DATA = 12'b110011011110;
            14'b00_011001010110: DATA = 12'b110011011100;
            14'b00_011001010111: DATA = 12'b110011011001;
            14'b00_011001011000: DATA = 12'b110011010111;
            14'b00_011001011001: DATA = 12'b110011010100;
            14'b00_011001011010: DATA = 12'b110011010010;
            14'b00_011001011011: DATA = 12'b110011001111;
            14'b00_011001011100: DATA = 12'b110011001101;
            14'b00_011001011101: DATA = 12'b110011001010;
            14'b00_011001011110: DATA = 12'b110011001000;
            14'b00_011001011111: DATA = 12'b110011000101;
            14'b00_011001100000: DATA = 12'b110011000011;
            14'b00_011001100001: DATA = 12'b110011000000;
            14'b00_011001100010: DATA = 12'b110010111110;
            14'b00_011001100011: DATA = 12'b110010111011;
            14'b00_011001100100: DATA = 12'b110010111001;
            14'b00_011001100101: DATA = 12'b110010110110;
            14'b00_011001100110: DATA = 12'b110010110100;
            14'b00_011001100111: DATA = 12'b110010110001;
            14'b00_011001101000: DATA = 12'b110010101111;
            14'b00_011001101001: DATA = 12'b110010101100;
            14'b00_011001101010: DATA = 12'b110010101010;
            14'b00_011001101011: DATA = 12'b110010100111;
            14'b00_011001101100: DATA = 12'b110010100100;
            14'b00_011001101101: DATA = 12'b110010100010;
            14'b00_011001101110: DATA = 12'b110010011111;
            14'b00_011001101111: DATA = 12'b110010011101;
            14'b00_011001110000: DATA = 12'b110010011010;
            14'b00_011001110001: DATA = 12'b110010011000;
            14'b00_011001110010: DATA = 12'b110010010101;
            14'b00_011001110011: DATA = 12'b110010010010;
            14'b00_011001110100: DATA = 12'b110010010000;
            14'b00_011001110101: DATA = 12'b110010001101;
            14'b00_011001110110: DATA = 12'b110010001011;
            14'b00_011001110111: DATA = 12'b110010001000;
            14'b00_011001111000: DATA = 12'b110010000110;
            14'b00_011001111001: DATA = 12'b110010000011;
            14'b00_011001111010: DATA = 12'b110010000000;
            14'b00_011001111011: DATA = 12'b110001111110;
            14'b00_011001111100: DATA = 12'b110001111011;
            14'b00_011001111101: DATA = 12'b110001111001;
            14'b00_011001111110: DATA = 12'b110001110110;
            14'b00_011001111111: DATA = 12'b110001110011;
            14'b00_011010000000: DATA = 12'b110001110001;
            14'b00_011010000001: DATA = 12'b110001101110;
            14'b00_011010000010: DATA = 12'b110001101100;
            14'b00_011010000011: DATA = 12'b110001101001;
            14'b00_011010000100: DATA = 12'b110001100110;
            14'b00_011010000101: DATA = 12'b110001100100;
            14'b00_011010000110: DATA = 12'b110001100001;
            14'b00_011010000111: DATA = 12'b110001011110;
            14'b00_011010001000: DATA = 12'b110001011100;
            14'b00_011010001001: DATA = 12'b110001011001;
            14'b00_011010001010: DATA = 12'b110001010111;
            14'b00_011010001011: DATA = 12'b110001010100;
            14'b00_011010001100: DATA = 12'b110001010001;
            14'b00_011010001101: DATA = 12'b110001001111;
            14'b00_011010001110: DATA = 12'b110001001100;
            14'b00_011010001111: DATA = 12'b110001001001;
            14'b00_011010010000: DATA = 12'b110001000111;
            14'b00_011010010001: DATA = 12'b110001000100;
            14'b00_011010010010: DATA = 12'b110001000001;
            14'b00_011010010011: DATA = 12'b110000111111;
            14'b00_011010010100: DATA = 12'b110000111100;
            14'b00_011010010101: DATA = 12'b110000111001;
            14'b00_011010010110: DATA = 12'b110000110111;
            14'b00_011010010111: DATA = 12'b110000110100;
            14'b00_011010011000: DATA = 12'b110000110001;
            14'b00_011010011001: DATA = 12'b110000101111;
            14'b00_011010011010: DATA = 12'b110000101100;
            14'b00_011010011011: DATA = 12'b110000101001;
            14'b00_011010011100: DATA = 12'b110000100111;
            14'b00_011010011101: DATA = 12'b110000100100;
            14'b00_011010011110: DATA = 12'b110000100001;
            14'b00_011010011111: DATA = 12'b110000011111;
            14'b00_011010100000: DATA = 12'b110000011100;
            14'b00_011010100001: DATA = 12'b110000011001;
            14'b00_011010100010: DATA = 12'b110000010110;
            14'b00_011010100011: DATA = 12'b110000010100;
            14'b00_011010100100: DATA = 12'b110000010001;
            14'b00_011010100101: DATA = 12'b110000001110;
            14'b00_011010100110: DATA = 12'b110000001100;
            14'b00_011010100111: DATA = 12'b110000001001;
            14'b00_011010101000: DATA = 12'b110000000110;
            14'b00_011010101001: DATA = 12'b110000000100;
            14'b00_011010101010: DATA = 12'b110000000001;
            14'b00_011010101011: DATA = 12'b101111111110;
            14'b00_011010101100: DATA = 12'b101111111011;
            14'b00_011010101101: DATA = 12'b101111111001;
            14'b00_011010101110: DATA = 12'b101111110110;
            14'b00_011010101111: DATA = 12'b101111110011;
            14'b00_011010110000: DATA = 12'b101111110000;
            14'b00_011010110001: DATA = 12'b101111101110;
            14'b00_011010110010: DATA = 12'b101111101011;
            14'b00_011010110011: DATA = 12'b101111101000;
            14'b00_011010110100: DATA = 12'b101111100110;
            14'b00_011010110101: DATA = 12'b101111100011;
            14'b00_011010110110: DATA = 12'b101111100000;
            14'b00_011010110111: DATA = 12'b101111011101;
            14'b00_011010111000: DATA = 12'b101111011011;
            14'b00_011010111001: DATA = 12'b101111011000;
            14'b00_011010111010: DATA = 12'b101111010101;
            14'b00_011010111011: DATA = 12'b101111010010;
            14'b00_011010111100: DATA = 12'b101111010000;
            14'b00_011010111101: DATA = 12'b101111001101;
            14'b00_011010111110: DATA = 12'b101111001010;
            14'b00_011010111111: DATA = 12'b101111000111;
            14'b00_011011000000: DATA = 12'b101111000100;
            14'b00_011011000001: DATA = 12'b101111000010;
            14'b00_011011000010: DATA = 12'b101110111111;
            14'b00_011011000011: DATA = 12'b101110111100;
            14'b00_011011000100: DATA = 12'b101110111001;
            14'b00_011011000101: DATA = 12'b101110110111;
            14'b00_011011000110: DATA = 12'b101110110100;
            14'b00_011011000111: DATA = 12'b101110110001;
            14'b00_011011001000: DATA = 12'b101110101110;
            14'b00_011011001001: DATA = 12'b101110101011;
            14'b00_011011001010: DATA = 12'b101110101001;
            14'b00_011011001011: DATA = 12'b101110100110;
            14'b00_011011001100: DATA = 12'b101110100011;
            14'b00_011011001101: DATA = 12'b101110100000;
            14'b00_011011001110: DATA = 12'b101110011101;
            14'b00_011011001111: DATA = 12'b101110011011;
            14'b00_011011010000: DATA = 12'b101110011000;
            14'b00_011011010001: DATA = 12'b101110010101;
            14'b00_011011010010: DATA = 12'b101110010010;
            14'b00_011011010011: DATA = 12'b101110001111;
            14'b00_011011010100: DATA = 12'b101110001101;
            14'b00_011011010101: DATA = 12'b101110001010;
            14'b00_011011010110: DATA = 12'b101110000111;
            14'b00_011011010111: DATA = 12'b101110000100;
            14'b00_011011011000: DATA = 12'b101110000001;
            14'b00_011011011001: DATA = 12'b101101111111;
            14'b00_011011011010: DATA = 12'b101101111100;
            14'b00_011011011011: DATA = 12'b101101111001;
            14'b00_011011011100: DATA = 12'b101101110110;
            14'b00_011011011101: DATA = 12'b101101110011;
            14'b00_011011011110: DATA = 12'b101101110000;
            14'b00_011011011111: DATA = 12'b101101101110;
            14'b00_011011100000: DATA = 12'b101101101011;
            14'b00_011011100001: DATA = 12'b101101101000;
            14'b00_011011100010: DATA = 12'b101101100101;
            14'b00_011011100011: DATA = 12'b101101100010;
            14'b00_011011100100: DATA = 12'b101101011111;
            14'b00_011011100101: DATA = 12'b101101011100;
            14'b00_011011100110: DATA = 12'b101101011010;
            14'b00_011011100111: DATA = 12'b101101010111;
            14'b00_011011101000: DATA = 12'b101101010100;
            14'b00_011011101001: DATA = 12'b101101010001;
            14'b00_011011101010: DATA = 12'b101101001110;
            14'b00_011011101011: DATA = 12'b101101001011;
            14'b00_011011101100: DATA = 12'b101101001000;
            14'b00_011011101101: DATA = 12'b101101000110;
            14'b00_011011101110: DATA = 12'b101101000011;
            14'b00_011011101111: DATA = 12'b101101000000;
            14'b00_011011110000: DATA = 12'b101100111101;
            14'b00_011011110001: DATA = 12'b101100111010;
            14'b00_011011110010: DATA = 12'b101100110111;
            14'b00_011011110011: DATA = 12'b101100110100;
            14'b00_011011110100: DATA = 12'b101100110010;
            14'b00_011011110101: DATA = 12'b101100101111;
            14'b00_011011110110: DATA = 12'b101100101100;
            14'b00_011011110111: DATA = 12'b101100101001;
            14'b00_011011111000: DATA = 12'b101100100110;
            14'b00_011011111001: DATA = 12'b101100100011;
            14'b00_011011111010: DATA = 12'b101100100000;
            14'b00_011011111011: DATA = 12'b101100011101;
            14'b00_011011111100: DATA = 12'b101100011010;
            14'b00_011011111101: DATA = 12'b101100011000;
            14'b00_011011111110: DATA = 12'b101100010101;
            14'b00_011011111111: DATA = 12'b101100010010;
            14'b00_011100000000: DATA = 12'b101100001111;
            14'b00_011100000001: DATA = 12'b101100001100;
            14'b00_011100000010: DATA = 12'b101100001001;
            14'b00_011100000011: DATA = 12'b101100000110;
            14'b00_011100000100: DATA = 12'b101100000011;
            14'b00_011100000101: DATA = 12'b101100000000;
            14'b00_011100000110: DATA = 12'b101011111101;
            14'b00_011100000111: DATA = 12'b101011111011;
            14'b00_011100001000: DATA = 12'b101011111000;
            14'b00_011100001001: DATA = 12'b101011110101;
            14'b00_011100001010: DATA = 12'b101011110010;
            14'b00_011100001011: DATA = 12'b101011101111;
            14'b00_011100001100: DATA = 12'b101011101100;
            14'b00_011100001101: DATA = 12'b101011101001;
            14'b00_011100001110: DATA = 12'b101011100110;
            14'b00_011100001111: DATA = 12'b101011100011;
            14'b00_011100010000: DATA = 12'b101011100000;
            14'b00_011100010001: DATA = 12'b101011011101;
            14'b00_011100010010: DATA = 12'b101011011010;
            14'b00_011100010011: DATA = 12'b101011010111;
            14'b00_011100010100: DATA = 12'b101011010100;
            14'b00_011100010101: DATA = 12'b101011010010;
            14'b00_011100010110: DATA = 12'b101011001111;
            14'b00_011100010111: DATA = 12'b101011001100;
            14'b00_011100011000: DATA = 12'b101011001001;
            14'b00_011100011001: DATA = 12'b101011000110;
            14'b00_011100011010: DATA = 12'b101011000011;
            14'b00_011100011011: DATA = 12'b101011000000;
            14'b00_011100011100: DATA = 12'b101010111101;
            14'b00_011100011101: DATA = 12'b101010111010;
            14'b00_011100011110: DATA = 12'b101010110111;
            14'b00_011100011111: DATA = 12'b101010110100;
            14'b00_011100100000: DATA = 12'b101010110001;
            14'b00_011100100001: DATA = 12'b101010101110;
            14'b00_011100100010: DATA = 12'b101010101011;
            14'b00_011100100011: DATA = 12'b101010101000;
            14'b00_011100100100: DATA = 12'b101010100101;
            14'b00_011100100101: DATA = 12'b101010100010;
            14'b00_011100100110: DATA = 12'b101010011111;
            14'b00_011100100111: DATA = 12'b101010011100;
            14'b00_011100101000: DATA = 12'b101010011001;
            14'b00_011100101001: DATA = 12'b101010010110;
            14'b00_011100101010: DATA = 12'b101010010011;
            14'b00_011100101011: DATA = 12'b101010010000;
            14'b00_011100101100: DATA = 12'b101010001110;
            14'b00_011100101101: DATA = 12'b101010001011;
            14'b00_011100101110: DATA = 12'b101010001000;
            14'b00_011100101111: DATA = 12'b101010000101;
            14'b00_011100110000: DATA = 12'b101010000010;
            14'b00_011100110001: DATA = 12'b101001111111;
            14'b00_011100110010: DATA = 12'b101001111100;
            14'b00_011100110011: DATA = 12'b101001111001;
            14'b00_011100110100: DATA = 12'b101001110110;
            14'b00_011100110101: DATA = 12'b101001110011;
            14'b00_011100110110: DATA = 12'b101001110000;
            14'b00_011100110111: DATA = 12'b101001101101;
            14'b00_011100111000: DATA = 12'b101001101010;
            14'b00_011100111001: DATA = 12'b101001100111;
            14'b00_011100111010: DATA = 12'b101001100100;
            14'b00_011100111011: DATA = 12'b101001100001;
            14'b00_011100111100: DATA = 12'b101001011110;
            14'b00_011100111101: DATA = 12'b101001011011;
            14'b00_011100111110: DATA = 12'b101001011000;
            14'b00_011100111111: DATA = 12'b101001010101;
            14'b00_011101000000: DATA = 12'b101001010010;
            14'b00_011101000001: DATA = 12'b101001001111;
            14'b00_011101000010: DATA = 12'b101001001100;
            14'b00_011101000011: DATA = 12'b101001001001;
            14'b00_011101000100: DATA = 12'b101001000110;
            14'b00_011101000101: DATA = 12'b101001000011;
            14'b00_011101000110: DATA = 12'b101001000000;
            14'b00_011101000111: DATA = 12'b101000111101;
            14'b00_011101001000: DATA = 12'b101000111010;
            14'b00_011101001001: DATA = 12'b101000110111;
            14'b00_011101001010: DATA = 12'b101000110100;
            14'b00_011101001011: DATA = 12'b101000110001;
            14'b00_011101001100: DATA = 12'b101000101110;
            14'b00_011101001101: DATA = 12'b101000101011;
            14'b00_011101001110: DATA = 12'b101000101000;
            14'b00_011101001111: DATA = 12'b101000100100;
            14'b00_011101010000: DATA = 12'b101000100001;
            14'b00_011101010001: DATA = 12'b101000011110;
            14'b00_011101010010: DATA = 12'b101000011011;
            14'b00_011101010011: DATA = 12'b101000011000;
            14'b00_011101010100: DATA = 12'b101000010101;
            14'b00_011101010101: DATA = 12'b101000010010;
            14'b00_011101010110: DATA = 12'b101000001111;
            14'b00_011101010111: DATA = 12'b101000001100;
            14'b00_011101011000: DATA = 12'b101000001001;
            14'b00_011101011001: DATA = 12'b101000000110;
            14'b00_011101011010: DATA = 12'b101000000011;
            14'b00_011101011011: DATA = 12'b101000000000;
            14'b00_011101011100: DATA = 12'b100111111101;
            14'b00_011101011101: DATA = 12'b100111111010;
            14'b00_011101011110: DATA = 12'b100111110111;
            14'b00_011101011111: DATA = 12'b100111110100;
            14'b00_011101100000: DATA = 12'b100111110001;
            14'b00_011101100001: DATA = 12'b100111101110;
            14'b00_011101100010: DATA = 12'b100111101011;
            14'b00_011101100011: DATA = 12'b100111101000;
            14'b00_011101100100: DATA = 12'b100111100101;
            14'b00_011101100101: DATA = 12'b100111100010;
            14'b00_011101100110: DATA = 12'b100111011111;
            14'b00_011101100111: DATA = 12'b100111011100;
            14'b00_011101101000: DATA = 12'b100111011000;
            14'b00_011101101001: DATA = 12'b100111010101;
            14'b00_011101101010: DATA = 12'b100111010010;
            14'b00_011101101011: DATA = 12'b100111001111;
            14'b00_011101101100: DATA = 12'b100111001100;
            14'b00_011101101101: DATA = 12'b100111001001;
            14'b00_011101101110: DATA = 12'b100111000110;
            14'b00_011101101111: DATA = 12'b100111000011;
            14'b00_011101110000: DATA = 12'b100111000000;
            14'b00_011101110001: DATA = 12'b100110111101;
            14'b00_011101110010: DATA = 12'b100110111010;
            14'b00_011101110011: DATA = 12'b100110110111;
            14'b00_011101110100: DATA = 12'b100110110100;
            14'b00_011101110101: DATA = 12'b100110110001;
            14'b00_011101110110: DATA = 12'b100110101110;
            14'b00_011101110111: DATA = 12'b100110101011;
            14'b00_011101111000: DATA = 12'b100110100111;
            14'b00_011101111001: DATA = 12'b100110100100;
            14'b00_011101111010: DATA = 12'b100110100001;
            14'b00_011101111011: DATA = 12'b100110011110;
            14'b00_011101111100: DATA = 12'b100110011011;
            14'b00_011101111101: DATA = 12'b100110011000;
            14'b00_011101111110: DATA = 12'b100110010101;
            14'b00_011101111111: DATA = 12'b100110010010;
            14'b00_011110000000: DATA = 12'b100110001111;
            14'b00_011110000001: DATA = 12'b100110001100;
            14'b00_011110000010: DATA = 12'b100110001001;
            14'b00_011110000011: DATA = 12'b100110000110;
            14'b00_011110000100: DATA = 12'b100110000011;
            14'b00_011110000101: DATA = 12'b100101111111;
            14'b00_011110000110: DATA = 12'b100101111100;
            14'b00_011110000111: DATA = 12'b100101111001;
            14'b00_011110001000: DATA = 12'b100101110110;
            14'b00_011110001001: DATA = 12'b100101110011;
            14'b00_011110001010: DATA = 12'b100101110000;
            14'b00_011110001011: DATA = 12'b100101101101;
            14'b00_011110001100: DATA = 12'b100101101010;
            14'b00_011110001101: DATA = 12'b100101100111;
            14'b00_011110001110: DATA = 12'b100101100100;
            14'b00_011110001111: DATA = 12'b100101100001;
            14'b00_011110010000: DATA = 12'b100101011101;
            14'b00_011110010001: DATA = 12'b100101011010;
            14'b00_011110010010: DATA = 12'b100101010111;
            14'b00_011110010011: DATA = 12'b100101010100;
            14'b00_011110010100: DATA = 12'b100101010001;
            14'b00_011110010101: DATA = 12'b100101001110;
            14'b00_011110010110: DATA = 12'b100101001011;
            14'b00_011110010111: DATA = 12'b100101001000;
            14'b00_011110011000: DATA = 12'b100101000101;
            14'b00_011110011001: DATA = 12'b100101000010;
            14'b00_011110011010: DATA = 12'b100100111110;
            14'b00_011110011011: DATA = 12'b100100111011;
            14'b00_011110011100: DATA = 12'b100100111000;
            14'b00_011110011101: DATA = 12'b100100110101;
            14'b00_011110011110: DATA = 12'b100100110010;
            14'b00_011110011111: DATA = 12'b100100101111;
            14'b00_011110100000: DATA = 12'b100100101100;
            14'b00_011110100001: DATA = 12'b100100101001;
            14'b00_011110100010: DATA = 12'b100100100110;
            14'b00_011110100011: DATA = 12'b100100100011;
            14'b00_011110100100: DATA = 12'b100100011111;
            14'b00_011110100101: DATA = 12'b100100011100;
            14'b00_011110100110: DATA = 12'b100100011001;
            14'b00_011110100111: DATA = 12'b100100010110;
            14'b00_011110101000: DATA = 12'b100100010011;
            14'b00_011110101001: DATA = 12'b100100010000;
            14'b00_011110101010: DATA = 12'b100100001101;
            14'b00_011110101011: DATA = 12'b100100001010;
            14'b00_011110101100: DATA = 12'b100100000111;
            14'b00_011110101101: DATA = 12'b100100000011;
            14'b00_011110101110: DATA = 12'b100100000000;
            14'b00_011110101111: DATA = 12'b100011111101;
            14'b00_011110110000: DATA = 12'b100011111010;
            14'b00_011110110001: DATA = 12'b100011110111;
            14'b00_011110110010: DATA = 12'b100011110100;
            14'b00_011110110011: DATA = 12'b100011110001;
            14'b00_011110110100: DATA = 12'b100011101110;
            14'b00_011110110101: DATA = 12'b100011101010;
            14'b00_011110110110: DATA = 12'b100011100111;
            14'b00_011110110111: DATA = 12'b100011100100;
            14'b00_011110111000: DATA = 12'b100011100001;
            14'b00_011110111001: DATA = 12'b100011011110;
            14'b00_011110111010: DATA = 12'b100011011011;
            14'b00_011110111011: DATA = 12'b100011011000;
            14'b00_011110111100: DATA = 12'b100011010101;
            14'b00_011110111101: DATA = 12'b100011010010;
            14'b00_011110111110: DATA = 12'b100011001110;
            14'b00_011110111111: DATA = 12'b100011001011;
            14'b00_011111000000: DATA = 12'b100011001000;
            14'b00_011111000001: DATA = 12'b100011000101;
            14'b00_011111000010: DATA = 12'b100011000010;
            14'b00_011111000011: DATA = 12'b100010111111;
            14'b00_011111000100: DATA = 12'b100010111100;
            14'b00_011111000101: DATA = 12'b100010111001;
            14'b00_011111000110: DATA = 12'b100010110101;
            14'b00_011111000111: DATA = 12'b100010110010;
            14'b00_011111001000: DATA = 12'b100010101111;
            14'b00_011111001001: DATA = 12'b100010101100;
            14'b00_011111001010: DATA = 12'b100010101001;
            14'b00_011111001011: DATA = 12'b100010100110;
            14'b00_011111001100: DATA = 12'b100010100011;
            14'b00_011111001101: DATA = 12'b100010011111;
            14'b00_011111001110: DATA = 12'b100010011100;
            14'b00_011111001111: DATA = 12'b100010011001;
            14'b00_011111010000: DATA = 12'b100010010110;
            14'b00_011111010001: DATA = 12'b100010010011;
            14'b00_011111010010: DATA = 12'b100010010000;
            14'b00_011111010011: DATA = 12'b100010001101;
            14'b00_011111010100: DATA = 12'b100010001010;
            14'b00_011111010101: DATA = 12'b100010000110;
            14'b00_011111010110: DATA = 12'b100010000011;
            14'b00_011111010111: DATA = 12'b100010000000;
            14'b00_011111011000: DATA = 12'b100001111101;
            14'b00_011111011001: DATA = 12'b100001111010;
            14'b00_011111011010: DATA = 12'b100001110111;
            14'b00_011111011011: DATA = 12'b100001110100;
            14'b00_011111011100: DATA = 12'b100001110000;
            14'b00_011111011101: DATA = 12'b100001101101;
            14'b00_011111011110: DATA = 12'b100001101010;
            14'b00_011111011111: DATA = 12'b100001100111;
            14'b00_011111100000: DATA = 12'b100001100100;
            14'b00_011111100001: DATA = 12'b100001100001;
            14'b00_011111100010: DATA = 12'b100001011110;
            14'b00_011111100011: DATA = 12'b100001011011;
            14'b00_011111100100: DATA = 12'b100001010111;
            14'b00_011111100101: DATA = 12'b100001010100;
            14'b00_011111100110: DATA = 12'b100001010001;
            14'b00_011111100111: DATA = 12'b100001001110;
            14'b00_011111101000: DATA = 12'b100001001011;
            14'b00_011111101001: DATA = 12'b100001001000;
            14'b00_011111101010: DATA = 12'b100001000101;
            14'b00_011111101011: DATA = 12'b100001000001;
            14'b00_011111101100: DATA = 12'b100000111110;
            14'b00_011111101101: DATA = 12'b100000111011;
            14'b00_011111101110: DATA = 12'b100000111000;
            14'b00_011111101111: DATA = 12'b100000110101;
            14'b00_011111110000: DATA = 12'b100000110010;
            14'b00_011111110001: DATA = 12'b100000101111;
            14'b00_011111110010: DATA = 12'b100000101011;
            14'b00_011111110011: DATA = 12'b100000101000;
            14'b00_011111110100: DATA = 12'b100000100101;
            14'b00_011111110101: DATA = 12'b100000100010;
            14'b00_011111110110: DATA = 12'b100000011111;
            14'b00_011111110111: DATA = 12'b100000011100;
            14'b00_011111111000: DATA = 12'b100000011001;
            14'b00_011111111001: DATA = 12'b100000010101;
            14'b00_011111111010: DATA = 12'b100000010010;
            14'b00_011111111011: DATA = 12'b100000001111;
            14'b00_011111111100: DATA = 12'b100000001100;
            14'b00_011111111101: DATA = 12'b100000001001;
            14'b00_011111111110: DATA = 12'b100000000110;
            14'b00_011111111111: DATA = 12'b100000000011;
            14'b00_100000000000: DATA = 12'b100000000000;
            14'b00_100000000001: DATA = 12'b011111111100;
            14'b00_100000000010: DATA = 12'b011111111001;
            14'b00_100000000011: DATA = 12'b011111110110;
            14'b00_100000000100: DATA = 12'b011111110011;
            14'b00_100000000101: DATA = 12'b011111110000;
            14'b00_100000000110: DATA = 12'b011111101101;
            14'b00_100000000111: DATA = 12'b011111101010;
            14'b00_100000001000: DATA = 12'b011111100110;
            14'b00_100000001001: DATA = 12'b011111100011;
            14'b00_100000001010: DATA = 12'b011111100000;
            14'b00_100000001011: DATA = 12'b011111011101;
            14'b00_100000001100: DATA = 12'b011111011010;
            14'b00_100000001101: DATA = 12'b011111010111;
            14'b00_100000001110: DATA = 12'b011111010100;
            14'b00_100000001111: DATA = 12'b011111010000;
            14'b00_100000010000: DATA = 12'b011111001101;
            14'b00_100000010001: DATA = 12'b011111001010;
            14'b00_100000010010: DATA = 12'b011111000111;
            14'b00_100000010011: DATA = 12'b011111000100;
            14'b00_100000010100: DATA = 12'b011111000001;
            14'b00_100000010101: DATA = 12'b011110111110;
            14'b00_100000010110: DATA = 12'b011110111010;
            14'b00_100000010111: DATA = 12'b011110110111;
            14'b00_100000011000: DATA = 12'b011110110100;
            14'b00_100000011001: DATA = 12'b011110110001;
            14'b00_100000011010: DATA = 12'b011110101110;
            14'b00_100000011011: DATA = 12'b011110101011;
            14'b00_100000011100: DATA = 12'b011110101000;
            14'b00_100000011101: DATA = 12'b011110100100;
            14'b00_100000011110: DATA = 12'b011110100001;
            14'b00_100000011111: DATA = 12'b011110011110;
            14'b00_100000100000: DATA = 12'b011110011011;
            14'b00_100000100001: DATA = 12'b011110011000;
            14'b00_100000100010: DATA = 12'b011110010101;
            14'b00_100000100011: DATA = 12'b011110010010;
            14'b00_100000100100: DATA = 12'b011110001111;
            14'b00_100000100101: DATA = 12'b011110001011;
            14'b00_100000100110: DATA = 12'b011110001000;
            14'b00_100000100111: DATA = 12'b011110000101;
            14'b00_100000101000: DATA = 12'b011110000010;
            14'b00_100000101001: DATA = 12'b011101111111;
            14'b00_100000101010: DATA = 12'b011101111100;
            14'b00_100000101011: DATA = 12'b011101111001;
            14'b00_100000101100: DATA = 12'b011101110101;
            14'b00_100000101101: DATA = 12'b011101110010;
            14'b00_100000101110: DATA = 12'b011101101111;
            14'b00_100000101111: DATA = 12'b011101101100;
            14'b00_100000110000: DATA = 12'b011101101001;
            14'b00_100000110001: DATA = 12'b011101100110;
            14'b00_100000110010: DATA = 12'b011101100011;
            14'b00_100000110011: DATA = 12'b011101100000;
            14'b00_100000110100: DATA = 12'b011101011100;
            14'b00_100000110101: DATA = 12'b011101011001;
            14'b00_100000110110: DATA = 12'b011101010110;
            14'b00_100000110111: DATA = 12'b011101010011;
            14'b00_100000111000: DATA = 12'b011101010000;
            14'b00_100000111001: DATA = 12'b011101001101;
            14'b00_100000111010: DATA = 12'b011101001010;
            14'b00_100000111011: DATA = 12'b011101000110;
            14'b00_100000111100: DATA = 12'b011101000011;
            14'b00_100000111101: DATA = 12'b011101000000;
            14'b00_100000111110: DATA = 12'b011100111101;
            14'b00_100000111111: DATA = 12'b011100111010;
            14'b00_100001000000: DATA = 12'b011100110111;
            14'b00_100001000001: DATA = 12'b011100110100;
            14'b00_100001000010: DATA = 12'b011100110001;
            14'b00_100001000011: DATA = 12'b011100101101;
            14'b00_100001000100: DATA = 12'b011100101010;
            14'b00_100001000101: DATA = 12'b011100100111;
            14'b00_100001000110: DATA = 12'b011100100100;
            14'b00_100001000111: DATA = 12'b011100100001;
            14'b00_100001001000: DATA = 12'b011100011110;
            14'b00_100001001001: DATA = 12'b011100011011;
            14'b00_100001001010: DATA = 12'b011100011000;
            14'b00_100001001011: DATA = 12'b011100010101;
            14'b00_100001001100: DATA = 12'b011100010001;
            14'b00_100001001101: DATA = 12'b011100001110;
            14'b00_100001001110: DATA = 12'b011100001011;
            14'b00_100001001111: DATA = 12'b011100001000;
            14'b00_100001010000: DATA = 12'b011100000101;
            14'b00_100001010001: DATA = 12'b011100000010;
            14'b00_100001010010: DATA = 12'b011011111111;
            14'b00_100001010011: DATA = 12'b011011111100;
            14'b00_100001010100: DATA = 12'b011011111000;
            14'b00_100001010101: DATA = 12'b011011110101;
            14'b00_100001010110: DATA = 12'b011011110010;
            14'b00_100001010111: DATA = 12'b011011101111;
            14'b00_100001011000: DATA = 12'b011011101100;
            14'b00_100001011001: DATA = 12'b011011101001;
            14'b00_100001011010: DATA = 12'b011011100110;
            14'b00_100001011011: DATA = 12'b011011100011;
            14'b00_100001011100: DATA = 12'b011011100000;
            14'b00_100001011101: DATA = 12'b011011011100;
            14'b00_100001011110: DATA = 12'b011011011001;
            14'b00_100001011111: DATA = 12'b011011010110;
            14'b00_100001100000: DATA = 12'b011011010011;
            14'b00_100001100001: DATA = 12'b011011010000;
            14'b00_100001100010: DATA = 12'b011011001101;
            14'b00_100001100011: DATA = 12'b011011001010;
            14'b00_100001100100: DATA = 12'b011011000111;
            14'b00_100001100101: DATA = 12'b011011000100;
            14'b00_100001100110: DATA = 12'b011011000001;
            14'b00_100001100111: DATA = 12'b011010111101;
            14'b00_100001101000: DATA = 12'b011010111010;
            14'b00_100001101001: DATA = 12'b011010110111;
            14'b00_100001101010: DATA = 12'b011010110100;
            14'b00_100001101011: DATA = 12'b011010110001;
            14'b00_100001101100: DATA = 12'b011010101110;
            14'b00_100001101101: DATA = 12'b011010101011;
            14'b00_100001101110: DATA = 12'b011010101000;
            14'b00_100001101111: DATA = 12'b011010100101;
            14'b00_100001110000: DATA = 12'b011010100010;
            14'b00_100001110001: DATA = 12'b011010011110;
            14'b00_100001110010: DATA = 12'b011010011011;
            14'b00_100001110011: DATA = 12'b011010011000;
            14'b00_100001110100: DATA = 12'b011010010101;
            14'b00_100001110101: DATA = 12'b011010010010;
            14'b00_100001110110: DATA = 12'b011010001111;
            14'b00_100001110111: DATA = 12'b011010001100;
            14'b00_100001111000: DATA = 12'b011010001001;
            14'b00_100001111001: DATA = 12'b011010000110;
            14'b00_100001111010: DATA = 12'b011010000011;
            14'b00_100001111011: DATA = 12'b011010000000;
            14'b00_100001111100: DATA = 12'b011001111100;
            14'b00_100001111101: DATA = 12'b011001111001;
            14'b00_100001111110: DATA = 12'b011001110110;
            14'b00_100001111111: DATA = 12'b011001110011;
            14'b00_100010000000: DATA = 12'b011001110000;
            14'b00_100010000001: DATA = 12'b011001101101;
            14'b00_100010000010: DATA = 12'b011001101010;
            14'b00_100010000011: DATA = 12'b011001100111;
            14'b00_100010000100: DATA = 12'b011001100100;
            14'b00_100010000101: DATA = 12'b011001100001;
            14'b00_100010000110: DATA = 12'b011001011110;
            14'b00_100010000111: DATA = 12'b011001011011;
            14'b00_100010001000: DATA = 12'b011001011000;
            14'b00_100010001001: DATA = 12'b011001010100;
            14'b00_100010001010: DATA = 12'b011001010001;
            14'b00_100010001011: DATA = 12'b011001001110;
            14'b00_100010001100: DATA = 12'b011001001011;
            14'b00_100010001101: DATA = 12'b011001001000;
            14'b00_100010001110: DATA = 12'b011001000101;
            14'b00_100010001111: DATA = 12'b011001000010;
            14'b00_100010010000: DATA = 12'b011000111111;
            14'b00_100010010001: DATA = 12'b011000111100;
            14'b00_100010010010: DATA = 12'b011000111001;
            14'b00_100010010011: DATA = 12'b011000110110;
            14'b00_100010010100: DATA = 12'b011000110011;
            14'b00_100010010101: DATA = 12'b011000110000;
            14'b00_100010010110: DATA = 12'b011000101101;
            14'b00_100010010111: DATA = 12'b011000101010;
            14'b00_100010011000: DATA = 12'b011000100111;
            14'b00_100010011001: DATA = 12'b011000100011;
            14'b00_100010011010: DATA = 12'b011000100000;
            14'b00_100010011011: DATA = 12'b011000011101;
            14'b00_100010011100: DATA = 12'b011000011010;
            14'b00_100010011101: DATA = 12'b011000010111;
            14'b00_100010011110: DATA = 12'b011000010100;
            14'b00_100010011111: DATA = 12'b011000010001;
            14'b00_100010100000: DATA = 12'b011000001110;
            14'b00_100010100001: DATA = 12'b011000001011;
            14'b00_100010100010: DATA = 12'b011000001000;
            14'b00_100010100011: DATA = 12'b011000000101;
            14'b00_100010100100: DATA = 12'b011000000010;
            14'b00_100010100101: DATA = 12'b010111111111;
            14'b00_100010100110: DATA = 12'b010111111100;
            14'b00_100010100111: DATA = 12'b010111111001;
            14'b00_100010101000: DATA = 12'b010111110110;
            14'b00_100010101001: DATA = 12'b010111110011;
            14'b00_100010101010: DATA = 12'b010111110000;
            14'b00_100010101011: DATA = 12'b010111101101;
            14'b00_100010101100: DATA = 12'b010111101010;
            14'b00_100010101101: DATA = 12'b010111100111;
            14'b00_100010101110: DATA = 12'b010111100100;
            14'b00_100010101111: DATA = 12'b010111100001;
            14'b00_100010110000: DATA = 12'b010111011110;
            14'b00_100010110001: DATA = 12'b010111011011;
            14'b00_100010110010: DATA = 12'b010111010111;
            14'b00_100010110011: DATA = 12'b010111010100;
            14'b00_100010110100: DATA = 12'b010111010001;
            14'b00_100010110101: DATA = 12'b010111001110;
            14'b00_100010110110: DATA = 12'b010111001011;
            14'b00_100010110111: DATA = 12'b010111001000;
            14'b00_100010111000: DATA = 12'b010111000101;
            14'b00_100010111001: DATA = 12'b010111000010;
            14'b00_100010111010: DATA = 12'b010110111111;
            14'b00_100010111011: DATA = 12'b010110111100;
            14'b00_100010111100: DATA = 12'b010110111001;
            14'b00_100010111101: DATA = 12'b010110110110;
            14'b00_100010111110: DATA = 12'b010110110011;
            14'b00_100010111111: DATA = 12'b010110110000;
            14'b00_100011000000: DATA = 12'b010110101101;
            14'b00_100011000001: DATA = 12'b010110101010;
            14'b00_100011000010: DATA = 12'b010110100111;
            14'b00_100011000011: DATA = 12'b010110100100;
            14'b00_100011000100: DATA = 12'b010110100001;
            14'b00_100011000101: DATA = 12'b010110011110;
            14'b00_100011000110: DATA = 12'b010110011011;
            14'b00_100011000111: DATA = 12'b010110011000;
            14'b00_100011001000: DATA = 12'b010110010101;
            14'b00_100011001001: DATA = 12'b010110010010;
            14'b00_100011001010: DATA = 12'b010110001111;
            14'b00_100011001011: DATA = 12'b010110001100;
            14'b00_100011001100: DATA = 12'b010110001001;
            14'b00_100011001101: DATA = 12'b010110000110;
            14'b00_100011001110: DATA = 12'b010110000011;
            14'b00_100011001111: DATA = 12'b010110000000;
            14'b00_100011010000: DATA = 12'b010101111101;
            14'b00_100011010001: DATA = 12'b010101111010;
            14'b00_100011010010: DATA = 12'b010101110111;
            14'b00_100011010011: DATA = 12'b010101110100;
            14'b00_100011010100: DATA = 12'b010101110001;
            14'b00_100011010101: DATA = 12'b010101101111;
            14'b00_100011010110: DATA = 12'b010101101100;
            14'b00_100011010111: DATA = 12'b010101101001;
            14'b00_100011011000: DATA = 12'b010101100110;
            14'b00_100011011001: DATA = 12'b010101100011;
            14'b00_100011011010: DATA = 12'b010101100000;
            14'b00_100011011011: DATA = 12'b010101011101;
            14'b00_100011011100: DATA = 12'b010101011010;
            14'b00_100011011101: DATA = 12'b010101010111;
            14'b00_100011011110: DATA = 12'b010101010100;
            14'b00_100011011111: DATA = 12'b010101010001;
            14'b00_100011100000: DATA = 12'b010101001110;
            14'b00_100011100001: DATA = 12'b010101001011;
            14'b00_100011100010: DATA = 12'b010101001000;
            14'b00_100011100011: DATA = 12'b010101000101;
            14'b00_100011100100: DATA = 12'b010101000010;
            14'b00_100011100101: DATA = 12'b010100111111;
            14'b00_100011100110: DATA = 12'b010100111100;
            14'b00_100011100111: DATA = 12'b010100111001;
            14'b00_100011101000: DATA = 12'b010100110110;
            14'b00_100011101001: DATA = 12'b010100110011;
            14'b00_100011101010: DATA = 12'b010100110000;
            14'b00_100011101011: DATA = 12'b010100101101;
            14'b00_100011101100: DATA = 12'b010100101011;
            14'b00_100011101101: DATA = 12'b010100101000;
            14'b00_100011101110: DATA = 12'b010100100101;
            14'b00_100011101111: DATA = 12'b010100100010;
            14'b00_100011110000: DATA = 12'b010100011111;
            14'b00_100011110001: DATA = 12'b010100011100;
            14'b00_100011110010: DATA = 12'b010100011001;
            14'b00_100011110011: DATA = 12'b010100010110;
            14'b00_100011110100: DATA = 12'b010100010011;
            14'b00_100011110101: DATA = 12'b010100010000;
            14'b00_100011110110: DATA = 12'b010100001101;
            14'b00_100011110111: DATA = 12'b010100001010;
            14'b00_100011111000: DATA = 12'b010100000111;
            14'b00_100011111001: DATA = 12'b010100000100;
            14'b00_100011111010: DATA = 12'b010100000010;
            14'b00_100011111011: DATA = 12'b010011111111;
            14'b00_100011111100: DATA = 12'b010011111100;
            14'b00_100011111101: DATA = 12'b010011111001;
            14'b00_100011111110: DATA = 12'b010011110110;
            14'b00_100011111111: DATA = 12'b010011110011;
            14'b00_100100000000: DATA = 12'b010011110000;
            14'b00_100100000001: DATA = 12'b010011101101;
            14'b00_100100000010: DATA = 12'b010011101010;
            14'b00_100100000011: DATA = 12'b010011100111;
            14'b00_100100000100: DATA = 12'b010011100101;
            14'b00_100100000101: DATA = 12'b010011100010;
            14'b00_100100000110: DATA = 12'b010011011111;
            14'b00_100100000111: DATA = 12'b010011011100;
            14'b00_100100001000: DATA = 12'b010011011001;
            14'b00_100100001001: DATA = 12'b010011010110;
            14'b00_100100001010: DATA = 12'b010011010011;
            14'b00_100100001011: DATA = 12'b010011010000;
            14'b00_100100001100: DATA = 12'b010011001101;
            14'b00_100100001101: DATA = 12'b010011001011;
            14'b00_100100001110: DATA = 12'b010011001000;
            14'b00_100100001111: DATA = 12'b010011000101;
            14'b00_100100010000: DATA = 12'b010011000010;
            14'b00_100100010001: DATA = 12'b010010111111;
            14'b00_100100010010: DATA = 12'b010010111100;
            14'b00_100100010011: DATA = 12'b010010111001;
            14'b00_100100010100: DATA = 12'b010010110111;
            14'b00_100100010101: DATA = 12'b010010110100;
            14'b00_100100010110: DATA = 12'b010010110001;
            14'b00_100100010111: DATA = 12'b010010101110;
            14'b00_100100011000: DATA = 12'b010010101011;
            14'b00_100100011001: DATA = 12'b010010101000;
            14'b00_100100011010: DATA = 12'b010010100101;
            14'b00_100100011011: DATA = 12'b010010100011;
            14'b00_100100011100: DATA = 12'b010010100000;
            14'b00_100100011101: DATA = 12'b010010011101;
            14'b00_100100011110: DATA = 12'b010010011010;
            14'b00_100100011111: DATA = 12'b010010010111;
            14'b00_100100100000: DATA = 12'b010010010100;
            14'b00_100100100001: DATA = 12'b010010010001;
            14'b00_100100100010: DATA = 12'b010010001111;
            14'b00_100100100011: DATA = 12'b010010001100;
            14'b00_100100100100: DATA = 12'b010010001001;
            14'b00_100100100101: DATA = 12'b010010000110;
            14'b00_100100100110: DATA = 12'b010010000011;
            14'b00_100100100111: DATA = 12'b010010000000;
            14'b00_100100101000: DATA = 12'b010001111110;
            14'b00_100100101001: DATA = 12'b010001111011;
            14'b00_100100101010: DATA = 12'b010001111000;
            14'b00_100100101011: DATA = 12'b010001110101;
            14'b00_100100101100: DATA = 12'b010001110010;
            14'b00_100100101101: DATA = 12'b010001110000;
            14'b00_100100101110: DATA = 12'b010001101101;
            14'b00_100100101111: DATA = 12'b010001101010;
            14'b00_100100110000: DATA = 12'b010001100111;
            14'b00_100100110001: DATA = 12'b010001100100;
            14'b00_100100110010: DATA = 12'b010001100010;
            14'b00_100100110011: DATA = 12'b010001011111;
            14'b00_100100110100: DATA = 12'b010001011100;
            14'b00_100100110101: DATA = 12'b010001011001;
            14'b00_100100110110: DATA = 12'b010001010110;
            14'b00_100100110111: DATA = 12'b010001010100;
            14'b00_100100111000: DATA = 12'b010001010001;
            14'b00_100100111001: DATA = 12'b010001001110;
            14'b00_100100111010: DATA = 12'b010001001011;
            14'b00_100100111011: DATA = 12'b010001001000;
            14'b00_100100111100: DATA = 12'b010001000110;
            14'b00_100100111101: DATA = 12'b010001000011;
            14'b00_100100111110: DATA = 12'b010001000000;
            14'b00_100100111111: DATA = 12'b010000111101;
            14'b00_100101000000: DATA = 12'b010000111011;
            14'b00_100101000001: DATA = 12'b010000111000;
            14'b00_100101000010: DATA = 12'b010000110101;
            14'b00_100101000011: DATA = 12'b010000110010;
            14'b00_100101000100: DATA = 12'b010000101111;
            14'b00_100101000101: DATA = 12'b010000101101;
            14'b00_100101000110: DATA = 12'b010000101010;
            14'b00_100101000111: DATA = 12'b010000100111;
            14'b00_100101001000: DATA = 12'b010000100100;
            14'b00_100101001001: DATA = 12'b010000100010;
            14'b00_100101001010: DATA = 12'b010000011111;
            14'b00_100101001011: DATA = 12'b010000011100;
            14'b00_100101001100: DATA = 12'b010000011001;
            14'b00_100101001101: DATA = 12'b010000010111;
            14'b00_100101001110: DATA = 12'b010000010100;
            14'b00_100101001111: DATA = 12'b010000010001;
            14'b00_100101010000: DATA = 12'b010000001111;
            14'b00_100101010001: DATA = 12'b010000001100;
            14'b00_100101010010: DATA = 12'b010000001001;
            14'b00_100101010011: DATA = 12'b010000000110;
            14'b00_100101010100: DATA = 12'b010000000100;
            14'b00_100101010101: DATA = 12'b010000000001;
            14'b00_100101010110: DATA = 12'b001111111110;
            14'b00_100101010111: DATA = 12'b001111111011;
            14'b00_100101011000: DATA = 12'b001111111001;
            14'b00_100101011001: DATA = 12'b001111110110;
            14'b00_100101011010: DATA = 12'b001111110011;
            14'b00_100101011011: DATA = 12'b001111110001;
            14'b00_100101011100: DATA = 12'b001111101110;
            14'b00_100101011101: DATA = 12'b001111101011;
            14'b00_100101011110: DATA = 12'b001111101001;
            14'b00_100101011111: DATA = 12'b001111100110;
            14'b00_100101100000: DATA = 12'b001111100011;
            14'b00_100101100001: DATA = 12'b001111100000;
            14'b00_100101100010: DATA = 12'b001111011110;
            14'b00_100101100011: DATA = 12'b001111011011;
            14'b00_100101100100: DATA = 12'b001111011000;
            14'b00_100101100101: DATA = 12'b001111010110;
            14'b00_100101100110: DATA = 12'b001111010011;
            14'b00_100101100111: DATA = 12'b001111010000;
            14'b00_100101101000: DATA = 12'b001111001110;
            14'b00_100101101001: DATA = 12'b001111001011;
            14'b00_100101101010: DATA = 12'b001111001000;
            14'b00_100101101011: DATA = 12'b001111000110;
            14'b00_100101101100: DATA = 12'b001111000011;
            14'b00_100101101101: DATA = 12'b001111000000;
            14'b00_100101101110: DATA = 12'b001110111110;
            14'b00_100101101111: DATA = 12'b001110111011;
            14'b00_100101110000: DATA = 12'b001110111000;
            14'b00_100101110001: DATA = 12'b001110110110;
            14'b00_100101110010: DATA = 12'b001110110011;
            14'b00_100101110011: DATA = 12'b001110110000;
            14'b00_100101110100: DATA = 12'b001110101110;
            14'b00_100101110101: DATA = 12'b001110101011;
            14'b00_100101110110: DATA = 12'b001110101000;
            14'b00_100101110111: DATA = 12'b001110100110;
            14'b00_100101111000: DATA = 12'b001110100011;
            14'b00_100101111001: DATA = 12'b001110100001;
            14'b00_100101111010: DATA = 12'b001110011110;
            14'b00_100101111011: DATA = 12'b001110011011;
            14'b00_100101111100: DATA = 12'b001110011001;
            14'b00_100101111101: DATA = 12'b001110010110;
            14'b00_100101111110: DATA = 12'b001110010011;
            14'b00_100101111111: DATA = 12'b001110010001;
            14'b00_100110000000: DATA = 12'b001110001110;
            14'b00_100110000001: DATA = 12'b001110001100;
            14'b00_100110000010: DATA = 12'b001110001001;
            14'b00_100110000011: DATA = 12'b001110000110;
            14'b00_100110000100: DATA = 12'b001110000100;
            14'b00_100110000101: DATA = 12'b001110000001;
            14'b00_100110000110: DATA = 12'b001101111111;
            14'b00_100110000111: DATA = 12'b001101111100;
            14'b00_100110001000: DATA = 12'b001101111001;
            14'b00_100110001001: DATA = 12'b001101110111;
            14'b00_100110001010: DATA = 12'b001101110100;
            14'b00_100110001011: DATA = 12'b001101110010;
            14'b00_100110001100: DATA = 12'b001101101111;
            14'b00_100110001101: DATA = 12'b001101101101;
            14'b00_100110001110: DATA = 12'b001101101010;
            14'b00_100110001111: DATA = 12'b001101100111;
            14'b00_100110010000: DATA = 12'b001101100101;
            14'b00_100110010001: DATA = 12'b001101100010;
            14'b00_100110010010: DATA = 12'b001101100000;
            14'b00_100110010011: DATA = 12'b001101011101;
            14'b00_100110010100: DATA = 12'b001101011011;
            14'b00_100110010101: DATA = 12'b001101011000;
            14'b00_100110010110: DATA = 12'b001101010101;
            14'b00_100110010111: DATA = 12'b001101010011;
            14'b00_100110011000: DATA = 12'b001101010000;
            14'b00_100110011001: DATA = 12'b001101001110;
            14'b00_100110011010: DATA = 12'b001101001011;
            14'b00_100110011011: DATA = 12'b001101001001;
            14'b00_100110011100: DATA = 12'b001101000110;
            14'b00_100110011101: DATA = 12'b001101000100;
            14'b00_100110011110: DATA = 12'b001101000001;
            14'b00_100110011111: DATA = 12'b001100111111;
            14'b00_100110100000: DATA = 12'b001100111100;
            14'b00_100110100001: DATA = 12'b001100111010;
            14'b00_100110100010: DATA = 12'b001100110111;
            14'b00_100110100011: DATA = 12'b001100110101;
            14'b00_100110100100: DATA = 12'b001100110010;
            14'b00_100110100101: DATA = 12'b001100110000;
            14'b00_100110100110: DATA = 12'b001100101101;
            14'b00_100110100111: DATA = 12'b001100101011;
            14'b00_100110101000: DATA = 12'b001100101000;
            14'b00_100110101001: DATA = 12'b001100100110;
            14'b00_100110101010: DATA = 12'b001100100011;
            14'b00_100110101011: DATA = 12'b001100100001;
            14'b00_100110101100: DATA = 12'b001100011110;
            14'b00_100110101101: DATA = 12'b001100011100;
            14'b00_100110101110: DATA = 12'b001100011001;
            14'b00_100110101111: DATA = 12'b001100010111;
            14'b00_100110110000: DATA = 12'b001100010100;
            14'b00_100110110001: DATA = 12'b001100010010;
            14'b00_100110110010: DATA = 12'b001100001111;
            14'b00_100110110011: DATA = 12'b001100001101;
            14'b00_100110110100: DATA = 12'b001100001010;
            14'b00_100110110101: DATA = 12'b001100001000;
            14'b00_100110110110: DATA = 12'b001100000101;
            14'b00_100110110111: DATA = 12'b001100000011;
            14'b00_100110111000: DATA = 12'b001100000000;
            14'b00_100110111001: DATA = 12'b001011111110;
            14'b00_100110111010: DATA = 12'b001011111100;
            14'b00_100110111011: DATA = 12'b001011111001;
            14'b00_100110111100: DATA = 12'b001011110111;
            14'b00_100110111101: DATA = 12'b001011110100;
            14'b00_100110111110: DATA = 12'b001011110010;
            14'b00_100110111111: DATA = 12'b001011101111;
            14'b00_100111000000: DATA = 12'b001011101101;
            14'b00_100111000001: DATA = 12'b001011101010;
            14'b00_100111000010: DATA = 12'b001011101000;
            14'b00_100111000011: DATA = 12'b001011100110;
            14'b00_100111000100: DATA = 12'b001011100011;
            14'b00_100111000101: DATA = 12'b001011100001;
            14'b00_100111000110: DATA = 12'b001011011110;
            14'b00_100111000111: DATA = 12'b001011011100;
            14'b00_100111001000: DATA = 12'b001011011010;
            14'b00_100111001001: DATA = 12'b001011010111;
            14'b00_100111001010: DATA = 12'b001011010101;
            14'b00_100111001011: DATA = 12'b001011010010;
            14'b00_100111001100: DATA = 12'b001011010000;
            14'b00_100111001101: DATA = 12'b001011001110;
            14'b00_100111001110: DATA = 12'b001011001011;
            14'b00_100111001111: DATA = 12'b001011001001;
            14'b00_100111010000: DATA = 12'b001011000110;
            14'b00_100111010001: DATA = 12'b001011000100;
            14'b00_100111010010: DATA = 12'b001011000010;
            14'b00_100111010011: DATA = 12'b001010111111;
            14'b00_100111010100: DATA = 12'b001010111101;
            14'b00_100111010101: DATA = 12'b001010111011;
            14'b00_100111010110: DATA = 12'b001010111000;
            14'b00_100111010111: DATA = 12'b001010110110;
            14'b00_100111011000: DATA = 12'b001010110100;
            14'b00_100111011001: DATA = 12'b001010110001;
            14'b00_100111011010: DATA = 12'b001010101111;
            14'b00_100111011011: DATA = 12'b001010101100;
            14'b00_100111011100: DATA = 12'b001010101010;
            14'b00_100111011101: DATA = 12'b001010101000;
            14'b00_100111011110: DATA = 12'b001010100101;
            14'b00_100111011111: DATA = 12'b001010100011;
            14'b00_100111100000: DATA = 12'b001010100001;
            14'b00_100111100001: DATA = 12'b001010011110;
            14'b00_100111100010: DATA = 12'b001010011100;
            14'b00_100111100011: DATA = 12'b001010011010;
            14'b00_100111100100: DATA = 12'b001010011000;
            14'b00_100111100101: DATA = 12'b001010010101;
            14'b00_100111100110: DATA = 12'b001010010011;
            14'b00_100111100111: DATA = 12'b001010010001;
            14'b00_100111101000: DATA = 12'b001010001110;
            14'b00_100111101001: DATA = 12'b001010001100;
            14'b00_100111101010: DATA = 12'b001010001010;
            14'b00_100111101011: DATA = 12'b001010000111;
            14'b00_100111101100: DATA = 12'b001010000101;
            14'b00_100111101101: DATA = 12'b001010000011;
            14'b00_100111101110: DATA = 12'b001010000001;
            14'b00_100111101111: DATA = 12'b001001111110;
            14'b00_100111110000: DATA = 12'b001001111100;
            14'b00_100111110001: DATA = 12'b001001111010;
            14'b00_100111110010: DATA = 12'b001001110111;
            14'b00_100111110011: DATA = 12'b001001110101;
            14'b00_100111110100: DATA = 12'b001001110011;
            14'b00_100111110101: DATA = 12'b001001110001;
            14'b00_100111110110: DATA = 12'b001001101110;
            14'b00_100111110111: DATA = 12'b001001101100;
            14'b00_100111111000: DATA = 12'b001001101010;
            14'b00_100111111001: DATA = 12'b001001101000;
            14'b00_100111111010: DATA = 12'b001001100101;
            14'b00_100111111011: DATA = 12'b001001100011;
            14'b00_100111111100: DATA = 12'b001001100001;
            14'b00_100111111101: DATA = 12'b001001011111;
            14'b00_100111111110: DATA = 12'b001001011100;
            14'b00_100111111111: DATA = 12'b001001011010;
            14'b00_101000000000: DATA = 12'b001001011000;
            14'b00_101000000001: DATA = 12'b001001010110;
            14'b00_101000000010: DATA = 12'b001001010100;
            14'b00_101000000011: DATA = 12'b001001010001;
            14'b00_101000000100: DATA = 12'b001001001111;
            14'b00_101000000101: DATA = 12'b001001001101;
            14'b00_101000000110: DATA = 12'b001001001011;
            14'b00_101000000111: DATA = 12'b001001001001;
            14'b00_101000001000: DATA = 12'b001001000110;
            14'b00_101000001001: DATA = 12'b001001000100;
            14'b00_101000001010: DATA = 12'b001001000010;
            14'b00_101000001011: DATA = 12'b001001000000;
            14'b00_101000001100: DATA = 12'b001000111110;
            14'b00_101000001101: DATA = 12'b001000111011;
            14'b00_101000001110: DATA = 12'b001000111001;
            14'b00_101000001111: DATA = 12'b001000110111;
            14'b00_101000010000: DATA = 12'b001000110101;
            14'b00_101000010001: DATA = 12'b001000110011;
            14'b00_101000010010: DATA = 12'b001000110001;
            14'b00_101000010011: DATA = 12'b001000101110;
            14'b00_101000010100: DATA = 12'b001000101100;
            14'b00_101000010101: DATA = 12'b001000101010;
            14'b00_101000010110: DATA = 12'b001000101000;
            14'b00_101000010111: DATA = 12'b001000100110;
            14'b00_101000011000: DATA = 12'b001000100100;
            14'b00_101000011001: DATA = 12'b001000100010;
            14'b00_101000011010: DATA = 12'b001000011111;
            14'b00_101000011011: DATA = 12'b001000011101;
            14'b00_101000011100: DATA = 12'b001000011011;
            14'b00_101000011101: DATA = 12'b001000011001;
            14'b00_101000011110: DATA = 12'b001000010111;
            14'b00_101000011111: DATA = 12'b001000010101;
            14'b00_101000100000: DATA = 12'b001000010011;
            14'b00_101000100001: DATA = 12'b001000010001;
            14'b00_101000100010: DATA = 12'b001000001111;
            14'b00_101000100011: DATA = 12'b001000001100;
            14'b00_101000100100: DATA = 12'b001000001010;
            14'b00_101000100101: DATA = 12'b001000001000;
            14'b00_101000100110: DATA = 12'b001000000110;
            14'b00_101000100111: DATA = 12'b001000000100;
            14'b00_101000101000: DATA = 12'b001000000010;
            14'b00_101000101001: DATA = 12'b001000000000;
            14'b00_101000101010: DATA = 12'b000111111110;
            14'b00_101000101011: DATA = 12'b000111111100;
            14'b00_101000101100: DATA = 12'b000111111010;
            14'b00_101000101101: DATA = 12'b000111111000;
            14'b00_101000101110: DATA = 12'b000111110110;
            14'b00_101000101111: DATA = 12'b000111110100;
            14'b00_101000110000: DATA = 12'b000111110001;
            14'b00_101000110001: DATA = 12'b000111101111;
            14'b00_101000110010: DATA = 12'b000111101101;
            14'b00_101000110011: DATA = 12'b000111101011;
            14'b00_101000110100: DATA = 12'b000111101001;
            14'b00_101000110101: DATA = 12'b000111100111;
            14'b00_101000110110: DATA = 12'b000111100101;
            14'b00_101000110111: DATA = 12'b000111100011;
            14'b00_101000111000: DATA = 12'b000111100001;
            14'b00_101000111001: DATA = 12'b000111011111;
            14'b00_101000111010: DATA = 12'b000111011101;
            14'b00_101000111011: DATA = 12'b000111011011;
            14'b00_101000111100: DATA = 12'b000111011001;
            14'b00_101000111101: DATA = 12'b000111010111;
            14'b00_101000111110: DATA = 12'b000111010101;
            14'b00_101000111111: DATA = 12'b000111010011;
            14'b00_101001000000: DATA = 12'b000111010001;
            14'b00_101001000001: DATA = 12'b000111001111;
            14'b00_101001000010: DATA = 12'b000111001101;
            14'b00_101001000011: DATA = 12'b000111001011;
            14'b00_101001000100: DATA = 12'b000111001001;
            14'b00_101001000101: DATA = 12'b000111000111;
            14'b00_101001000110: DATA = 12'b000111000101;
            14'b00_101001000111: DATA = 12'b000111000011;
            14'b00_101001001000: DATA = 12'b000111000001;
            14'b00_101001001001: DATA = 12'b000110111111;
            14'b00_101001001010: DATA = 12'b000110111101;
            14'b00_101001001011: DATA = 12'b000110111011;
            14'b00_101001001100: DATA = 12'b000110111010;
            14'b00_101001001101: DATA = 12'b000110111000;
            14'b00_101001001110: DATA = 12'b000110110110;
            14'b00_101001001111: DATA = 12'b000110110100;
            14'b00_101001010000: DATA = 12'b000110110010;
            14'b00_101001010001: DATA = 12'b000110110000;
            14'b00_101001010010: DATA = 12'b000110101110;
            14'b00_101001010011: DATA = 12'b000110101100;
            14'b00_101001010100: DATA = 12'b000110101010;
            14'b00_101001010101: DATA = 12'b000110101000;
            14'b00_101001010110: DATA = 12'b000110100110;
            14'b00_101001010111: DATA = 12'b000110100100;
            14'b00_101001011000: DATA = 12'b000110100010;
            14'b00_101001011001: DATA = 12'b000110100001;
            14'b00_101001011010: DATA = 12'b000110011111;
            14'b00_101001011011: DATA = 12'b000110011101;
            14'b00_101001011100: DATA = 12'b000110011011;
            14'b00_101001011101: DATA = 12'b000110011001;
            14'b00_101001011110: DATA = 12'b000110010111;
            14'b00_101001011111: DATA = 12'b000110010101;
            14'b00_101001100000: DATA = 12'b000110010011;
            14'b00_101001100001: DATA = 12'b000110010001;
            14'b00_101001100010: DATA = 12'b000110010000;
            14'b00_101001100011: DATA = 12'b000110001110;
            14'b00_101001100100: DATA = 12'b000110001100;
            14'b00_101001100101: DATA = 12'b000110001010;
            14'b00_101001100110: DATA = 12'b000110001000;
            14'b00_101001100111: DATA = 12'b000110000110;
            14'b00_101001101000: DATA = 12'b000110000100;
            14'b00_101001101001: DATA = 12'b000110000011;
            14'b00_101001101010: DATA = 12'b000110000001;
            14'b00_101001101011: DATA = 12'b000101111111;
            14'b00_101001101100: DATA = 12'b000101111101;
            14'b00_101001101101: DATA = 12'b000101111011;
            14'b00_101001101110: DATA = 12'b000101111010;
            14'b00_101001101111: DATA = 12'b000101111000;
            14'b00_101001110000: DATA = 12'b000101110110;
            14'b00_101001110001: DATA = 12'b000101110100;
            14'b00_101001110010: DATA = 12'b000101110010;
            14'b00_101001110011: DATA = 12'b000101110000;
            14'b00_101001110100: DATA = 12'b000101101111;
            14'b00_101001110101: DATA = 12'b000101101101;
            14'b00_101001110110: DATA = 12'b000101101011;
            14'b00_101001110111: DATA = 12'b000101101001;
            14'b00_101001111000: DATA = 12'b000101101000;
            14'b00_101001111001: DATA = 12'b000101100110;
            14'b00_101001111010: DATA = 12'b000101100100;
            14'b00_101001111011: DATA = 12'b000101100010;
            14'b00_101001111100: DATA = 12'b000101100000;
            14'b00_101001111101: DATA = 12'b000101011111;
            14'b00_101001111110: DATA = 12'b000101011101;
            14'b00_101001111111: DATA = 12'b000101011011;
            14'b00_101010000000: DATA = 12'b000101011001;
            14'b00_101010000001: DATA = 12'b000101011000;
            14'b00_101010000010: DATA = 12'b000101010110;
            14'b00_101010000011: DATA = 12'b000101010100;
            14'b00_101010000100: DATA = 12'b000101010011;
            14'b00_101010000101: DATA = 12'b000101010001;
            14'b00_101010000110: DATA = 12'b000101001111;
            14'b00_101010000111: DATA = 12'b000101001101;
            14'b00_101010001000: DATA = 12'b000101001100;
            14'b00_101010001001: DATA = 12'b000101001010;
            14'b00_101010001010: DATA = 12'b000101001000;
            14'b00_101010001011: DATA = 12'b000101000111;
            14'b00_101010001100: DATA = 12'b000101000101;
            14'b00_101010001101: DATA = 12'b000101000011;
            14'b00_101010001110: DATA = 12'b000101000001;
            14'b00_101010001111: DATA = 12'b000101000000;
            14'b00_101010010000: DATA = 12'b000100111110;
            14'b00_101010010001: DATA = 12'b000100111100;
            14'b00_101010010010: DATA = 12'b000100111011;
            14'b00_101010010011: DATA = 12'b000100111001;
            14'b00_101010010100: DATA = 12'b000100110111;
            14'b00_101010010101: DATA = 12'b000100110110;
            14'b00_101010010110: DATA = 12'b000100110100;
            14'b00_101010010111: DATA = 12'b000100110010;
            14'b00_101010011000: DATA = 12'b000100110001;
            14'b00_101010011001: DATA = 12'b000100101111;
            14'b00_101010011010: DATA = 12'b000100101101;
            14'b00_101010011011: DATA = 12'b000100101100;
            14'b00_101010011100: DATA = 12'b000100101010;
            14'b00_101010011101: DATA = 12'b000100101001;
            14'b00_101010011110: DATA = 12'b000100100111;
            14'b00_101010011111: DATA = 12'b000100100101;
            14'b00_101010100000: DATA = 12'b000100100100;
            14'b00_101010100001: DATA = 12'b000100100010;
            14'b00_101010100010: DATA = 12'b000100100001;
            14'b00_101010100011: DATA = 12'b000100011111;
            14'b00_101010100100: DATA = 12'b000100011101;
            14'b00_101010100101: DATA = 12'b000100011100;
            14'b00_101010100110: DATA = 12'b000100011010;
            14'b00_101010100111: DATA = 12'b000100011001;
            14'b00_101010101000: DATA = 12'b000100010111;
            14'b00_101010101001: DATA = 12'b000100010101;
            14'b00_101010101010: DATA = 12'b000100010100;
            14'b00_101010101011: DATA = 12'b000100010010;
            14'b00_101010101100: DATA = 12'b000100010001;
            14'b00_101010101101: DATA = 12'b000100001111;
            14'b00_101010101110: DATA = 12'b000100001110;
            14'b00_101010101111: DATA = 12'b000100001100;
            14'b00_101010110000: DATA = 12'b000100001010;
            14'b00_101010110001: DATA = 12'b000100001001;
            14'b00_101010110010: DATA = 12'b000100000111;
            14'b00_101010110011: DATA = 12'b000100000110;
            14'b00_101010110100: DATA = 12'b000100000100;
            14'b00_101010110101: DATA = 12'b000100000011;
            14'b00_101010110110: DATA = 12'b000100000001;
            14'b00_101010110111: DATA = 12'b000100000000;
            14'b00_101010111000: DATA = 12'b000011111110;
            14'b00_101010111001: DATA = 12'b000011111101;
            14'b00_101010111010: DATA = 12'b000011111011;
            14'b00_101010111011: DATA = 12'b000011111010;
            14'b00_101010111100: DATA = 12'b000011111000;
            14'b00_101010111101: DATA = 12'b000011110111;
            14'b00_101010111110: DATA = 12'b000011110101;
            14'b00_101010111111: DATA = 12'b000011110100;
            14'b00_101011000000: DATA = 12'b000011110010;
            14'b00_101011000001: DATA = 12'b000011110001;
            14'b00_101011000010: DATA = 12'b000011101111;
            14'b00_101011000011: DATA = 12'b000011101110;
            14'b00_101011000100: DATA = 12'b000011101100;
            14'b00_101011000101: DATA = 12'b000011101011;
            14'b00_101011000110: DATA = 12'b000011101001;
            14'b00_101011000111: DATA = 12'b000011101000;
            14'b00_101011001000: DATA = 12'b000011100111;
            14'b00_101011001001: DATA = 12'b000011100101;
            14'b00_101011001010: DATA = 12'b000011100100;
            14'b00_101011001011: DATA = 12'b000011100010;
            14'b00_101011001100: DATA = 12'b000011100001;
            14'b00_101011001101: DATA = 12'b000011011111;
            14'b00_101011001110: DATA = 12'b000011011110;
            14'b00_101011001111: DATA = 12'b000011011100;
            14'b00_101011010000: DATA = 12'b000011011011;
            14'b00_101011010001: DATA = 12'b000011011010;
            14'b00_101011010010: DATA = 12'b000011011000;
            14'b00_101011010011: DATA = 12'b000011010111;
            14'b00_101011010100: DATA = 12'b000011010101;
            14'b00_101011010101: DATA = 12'b000011010100;
            14'b00_101011010110: DATA = 12'b000011010011;
            14'b00_101011010111: DATA = 12'b000011010001;
            14'b00_101011011000: DATA = 12'b000011010000;
            14'b00_101011011001: DATA = 12'b000011001111;
            14'b00_101011011010: DATA = 12'b000011001101;
            14'b00_101011011011: DATA = 12'b000011001100;
            14'b00_101011011100: DATA = 12'b000011001010;
            14'b00_101011011101: DATA = 12'b000011001001;
            14'b00_101011011110: DATA = 12'b000011001000;
            14'b00_101011011111: DATA = 12'b000011000110;
            14'b00_101011100000: DATA = 12'b000011000101;
            14'b00_101011100001: DATA = 12'b000011000100;
            14'b00_101011100010: DATA = 12'b000011000010;
            14'b00_101011100011: DATA = 12'b000011000001;
            14'b00_101011100100: DATA = 12'b000011000000;
            14'b00_101011100101: DATA = 12'b000010111110;
            14'b00_101011100110: DATA = 12'b000010111101;
            14'b00_101011100111: DATA = 12'b000010111100;
            14'b00_101011101000: DATA = 12'b000010111010;
            14'b00_101011101001: DATA = 12'b000010111001;
            14'b00_101011101010: DATA = 12'b000010111000;
            14'b00_101011101011: DATA = 12'b000010110111;
            14'b00_101011101100: DATA = 12'b000010110101;
            14'b00_101011101101: DATA = 12'b000010110100;
            14'b00_101011101110: DATA = 12'b000010110011;
            14'b00_101011101111: DATA = 12'b000010110001;
            14'b00_101011110000: DATA = 12'b000010110000;
            14'b00_101011110001: DATA = 12'b000010101111;
            14'b00_101011110010: DATA = 12'b000010101110;
            14'b00_101011110011: DATA = 12'b000010101100;
            14'b00_101011110100: DATA = 12'b000010101011;
            14'b00_101011110101: DATA = 12'b000010101010;
            14'b00_101011110110: DATA = 12'b000010101001;
            14'b00_101011110111: DATA = 12'b000010100111;
            14'b00_101011111000: DATA = 12'b000010100110;
            14'b00_101011111001: DATA = 12'b000010100101;
            14'b00_101011111010: DATA = 12'b000010100100;
            14'b00_101011111011: DATA = 12'b000010100010;
            14'b00_101011111100: DATA = 12'b000010100001;
            14'b00_101011111101: DATA = 12'b000010100000;
            14'b00_101011111110: DATA = 12'b000010011111;
            14'b00_101011111111: DATA = 12'b000010011110;
            14'b00_101100000000: DATA = 12'b000010011100;
            14'b00_101100000001: DATA = 12'b000010011011;
            14'b00_101100000010: DATA = 12'b000010011010;
            14'b00_101100000011: DATA = 12'b000010011001;
            14'b00_101100000100: DATA = 12'b000010011000;
            14'b00_101100000101: DATA = 12'b000010010110;
            14'b00_101100000110: DATA = 12'b000010010101;
            14'b00_101100000111: DATA = 12'b000010010100;
            14'b00_101100001000: DATA = 12'b000010010011;
            14'b00_101100001001: DATA = 12'b000010010010;
            14'b00_101100001010: DATA = 12'b000010010001;
            14'b00_101100001011: DATA = 12'b000010001111;
            14'b00_101100001100: DATA = 12'b000010001110;
            14'b00_101100001101: DATA = 12'b000010001101;
            14'b00_101100001110: DATA = 12'b000010001100;
            14'b00_101100001111: DATA = 12'b000010001011;
            14'b00_101100010000: DATA = 12'b000010001010;
            14'b00_101100010001: DATA = 12'b000010001001;
            14'b00_101100010010: DATA = 12'b000010000111;
            14'b00_101100010011: DATA = 12'b000010000110;
            14'b00_101100010100: DATA = 12'b000010000101;
            14'b00_101100010101: DATA = 12'b000010000100;
            14'b00_101100010110: DATA = 12'b000010000011;
            14'b00_101100010111: DATA = 12'b000010000010;
            14'b00_101100011000: DATA = 12'b000010000001;
            14'b00_101100011001: DATA = 12'b000010000000;
            14'b00_101100011010: DATA = 12'b000001111111;
            14'b00_101100011011: DATA = 12'b000001111110;
            14'b00_101100011100: DATA = 12'b000001111100;
            14'b00_101100011101: DATA = 12'b000001111011;
            14'b00_101100011110: DATA = 12'b000001111010;
            14'b00_101100011111: DATA = 12'b000001111001;
            14'b00_101100100000: DATA = 12'b000001111000;
            14'b00_101100100001: DATA = 12'b000001110111;
            14'b00_101100100010: DATA = 12'b000001110110;
            14'b00_101100100011: DATA = 12'b000001110101;
            14'b00_101100100100: DATA = 12'b000001110100;
            14'b00_101100100101: DATA = 12'b000001110011;
            14'b00_101100100110: DATA = 12'b000001110010;
            14'b00_101100100111: DATA = 12'b000001110001;
            14'b00_101100101000: DATA = 12'b000001110000;
            14'b00_101100101001: DATA = 12'b000001101111;
            14'b00_101100101010: DATA = 12'b000001101110;
            14'b00_101100101011: DATA = 12'b000001101101;
            14'b00_101100101100: DATA = 12'b000001101100;
            14'b00_101100101101: DATA = 12'b000001101011;
            14'b00_101100101110: DATA = 12'b000001101010;
            14'b00_101100101111: DATA = 12'b000001101001;
            14'b00_101100110000: DATA = 12'b000001101000;
            14'b00_101100110001: DATA = 12'b000001100111;
            14'b00_101100110010: DATA = 12'b000001100110;
            14'b00_101100110011: DATA = 12'b000001100101;
            14'b00_101100110100: DATA = 12'b000001100100;
            14'b00_101100110101: DATA = 12'b000001100011;
            14'b00_101100110110: DATA = 12'b000001100010;
            14'b00_101100110111: DATA = 12'b000001100001;
            14'b00_101100111000: DATA = 12'b000001100000;
            14'b00_101100111001: DATA = 12'b000001011111;
            14'b00_101100111010: DATA = 12'b000001011110;
            14'b00_101100111011: DATA = 12'b000001011101;
            14'b00_101100111100: DATA = 12'b000001011100;
            14'b00_101100111101: DATA = 12'b000001011011;
            14'b00_101100111110: DATA = 12'b000001011010;
            14'b00_101100111111: DATA = 12'b000001011010;
            14'b00_101101000000: DATA = 12'b000001011001;
            14'b00_101101000001: DATA = 12'b000001011000;
            14'b00_101101000010: DATA = 12'b000001010111;
            14'b00_101101000011: DATA = 12'b000001010110;
            14'b00_101101000100: DATA = 12'b000001010101;
            14'b00_101101000101: DATA = 12'b000001010100;
            14'b00_101101000110: DATA = 12'b000001010011;
            14'b00_101101000111: DATA = 12'b000001010010;
            14'b00_101101001000: DATA = 12'b000001010001;
            14'b00_101101001001: DATA = 12'b000001010001;
            14'b00_101101001010: DATA = 12'b000001010000;
            14'b00_101101001011: DATA = 12'b000001001111;
            14'b00_101101001100: DATA = 12'b000001001110;
            14'b00_101101001101: DATA = 12'b000001001101;
            14'b00_101101001110: DATA = 12'b000001001100;
            14'b00_101101001111: DATA = 12'b000001001011;
            14'b00_101101010000: DATA = 12'b000001001011;
            14'b00_101101010001: DATA = 12'b000001001010;
            14'b00_101101010010: DATA = 12'b000001001001;
            14'b00_101101010011: DATA = 12'b000001001000;
            14'b00_101101010100: DATA = 12'b000001000111;
            14'b00_101101010101: DATA = 12'b000001000111;
            14'b00_101101010110: DATA = 12'b000001000110;
            14'b00_101101010111: DATA = 12'b000001000101;
            14'b00_101101011000: DATA = 12'b000001000100;
            14'b00_101101011001: DATA = 12'b000001000011;
            14'b00_101101011010: DATA = 12'b000001000011;
            14'b00_101101011011: DATA = 12'b000001000010;
            14'b00_101101011100: DATA = 12'b000001000001;
            14'b00_101101011101: DATA = 12'b000001000000;
            14'b00_101101011110: DATA = 12'b000000111111;
            14'b00_101101011111: DATA = 12'b000000111111;
            14'b00_101101100000: DATA = 12'b000000111110;
            14'b00_101101100001: DATA = 12'b000000111101;
            14'b00_101101100010: DATA = 12'b000000111100;
            14'b00_101101100011: DATA = 12'b000000111100;
            14'b00_101101100100: DATA = 12'b000000111011;
            14'b00_101101100101: DATA = 12'b000000111010;
            14'b00_101101100110: DATA = 12'b000000111001;
            14'b00_101101100111: DATA = 12'b000000111001;
            14'b00_101101101000: DATA = 12'b000000111000;
            14'b00_101101101001: DATA = 12'b000000110111;
            14'b00_101101101010: DATA = 12'b000000110110;
            14'b00_101101101011: DATA = 12'b000000110110;
            14'b00_101101101100: DATA = 12'b000000110101;
            14'b00_101101101101: DATA = 12'b000000110100;
            14'b00_101101101110: DATA = 12'b000000110100;
            14'b00_101101101111: DATA = 12'b000000110011;
            14'b00_101101110000: DATA = 12'b000000110010;
            14'b00_101101110001: DATA = 12'b000000110010;
            14'b00_101101110010: DATA = 12'b000000110001;
            14'b00_101101110011: DATA = 12'b000000110000;
            14'b00_101101110100: DATA = 12'b000000110000;
            14'b00_101101110101: DATA = 12'b000000101111;
            14'b00_101101110110: DATA = 12'b000000101110;
            14'b00_101101110111: DATA = 12'b000000101110;
            14'b00_101101111000: DATA = 12'b000000101101;
            14'b00_101101111001: DATA = 12'b000000101100;
            14'b00_101101111010: DATA = 12'b000000101100;
            14'b00_101101111011: DATA = 12'b000000101011;
            14'b00_101101111100: DATA = 12'b000000101010;
            14'b00_101101111101: DATA = 12'b000000101010;
            14'b00_101101111110: DATA = 12'b000000101001;
            14'b00_101101111111: DATA = 12'b000000101000;
            14'b00_101110000000: DATA = 12'b000000101000;
            14'b00_101110000001: DATA = 12'b000000100111;
            14'b00_101110000010: DATA = 12'b000000100111;
            14'b00_101110000011: DATA = 12'b000000100110;
            14'b00_101110000100: DATA = 12'b000000100101;
            14'b00_101110000101: DATA = 12'b000000100101;
            14'b00_101110000110: DATA = 12'b000000100100;
            14'b00_101110000111: DATA = 12'b000000100100;
            14'b00_101110001000: DATA = 12'b000000100011;
            14'b00_101110001001: DATA = 12'b000000100011;
            14'b00_101110001010: DATA = 12'b000000100010;
            14'b00_101110001011: DATA = 12'b000000100001;
            14'b00_101110001100: DATA = 12'b000000100001;
            14'b00_101110001101: DATA = 12'b000000100000;
            14'b00_101110001110: DATA = 12'b000000100000;
            14'b00_101110001111: DATA = 12'b000000011111;
            14'b00_101110010000: DATA = 12'b000000011111;
            14'b00_101110010001: DATA = 12'b000000011110;
            14'b00_101110010010: DATA = 12'b000000011110;
            14'b00_101110010011: DATA = 12'b000000011101;
            14'b00_101110010100: DATA = 12'b000000011101;
            14'b00_101110010101: DATA = 12'b000000011100;
            14'b00_101110010110: DATA = 12'b000000011100;
            14'b00_101110010111: DATA = 12'b000000011011;
            14'b00_101110011000: DATA = 12'b000000011010;
            14'b00_101110011001: DATA = 12'b000000011010;
            14'b00_101110011010: DATA = 12'b000000011010;
            14'b00_101110011011: DATA = 12'b000000011001;
            14'b00_101110011100: DATA = 12'b000000011001;
            14'b00_101110011101: DATA = 12'b000000011000;
            14'b00_101110011110: DATA = 12'b000000011000;
            14'b00_101110011111: DATA = 12'b000000010111;
            14'b00_101110100000: DATA = 12'b000000010111;
            14'b00_101110100001: DATA = 12'b000000010110;
            14'b00_101110100010: DATA = 12'b000000010110;
            14'b00_101110100011: DATA = 12'b000000010101;
            14'b00_101110100100: DATA = 12'b000000010101;
            14'b00_101110100101: DATA = 12'b000000010100;
            14'b00_101110100110: DATA = 12'b000000010100;
            14'b00_101110100111: DATA = 12'b000000010100;
            14'b00_101110101000: DATA = 12'b000000010011;
            14'b00_101110101001: DATA = 12'b000000010011;
            14'b00_101110101010: DATA = 12'b000000010010;
            14'b00_101110101011: DATA = 12'b000000010010;
            14'b00_101110101100: DATA = 12'b000000010001;
            14'b00_101110101101: DATA = 12'b000000010001;
            14'b00_101110101110: DATA = 12'b000000010001;
            14'b00_101110101111: DATA = 12'b000000010000;
            14'b00_101110110000: DATA = 12'b000000010000;
            14'b00_101110110001: DATA = 12'b000000010000;
            14'b00_101110110010: DATA = 12'b000000001111;
            14'b00_101110110011: DATA = 12'b000000001111;
            14'b00_101110110100: DATA = 12'b000000001110;
            14'b00_101110110101: DATA = 12'b000000001110;
            14'b00_101110110110: DATA = 12'b000000001110;
            14'b00_101110110111: DATA = 12'b000000001101;
            14'b00_101110111000: DATA = 12'b000000001101;
            14'b00_101110111001: DATA = 12'b000000001101;
            14'b00_101110111010: DATA = 12'b000000001100;
            14'b00_101110111011: DATA = 12'b000000001100;
            14'b00_101110111100: DATA = 12'b000000001100;
            14'b00_101110111101: DATA = 12'b000000001011;
            14'b00_101110111110: DATA = 12'b000000001011;
            14'b00_101110111111: DATA = 12'b000000001011;
            14'b00_101111000000: DATA = 12'b000000001010;
            14'b00_101111000001: DATA = 12'b000000001010;
            14'b00_101111000010: DATA = 12'b000000001010;
            14'b00_101111000011: DATA = 12'b000000001001;
            14'b00_101111000100: DATA = 12'b000000001001;
            14'b00_101111000101: DATA = 12'b000000001001;
            14'b00_101111000110: DATA = 12'b000000001001;
            14'b00_101111000111: DATA = 12'b000000001000;
            14'b00_101111001000: DATA = 12'b000000001000;
            14'b00_101111001001: DATA = 12'b000000001000;
            14'b00_101111001010: DATA = 12'b000000001000;
            14'b00_101111001011: DATA = 12'b000000000111;
            14'b00_101111001100: DATA = 12'b000000000111;
            14'b00_101111001101: DATA = 12'b000000000111;
            14'b00_101111001110: DATA = 12'b000000000111;
            14'b00_101111001111: DATA = 12'b000000000110;
            14'b00_101111010000: DATA = 12'b000000000110;
            14'b00_101111010001: DATA = 12'b000000000110;
            14'b00_101111010010: DATA = 12'b000000000110;
            14'b00_101111010011: DATA = 12'b000000000101;
            14'b00_101111010100: DATA = 12'b000000000101;
            14'b00_101111010101: DATA = 12'b000000000101;
            14'b00_101111010110: DATA = 12'b000000000101;
            14'b00_101111010111: DATA = 12'b000000000101;
            14'b00_101111011000: DATA = 12'b000000000100;
            14'b00_101111011001: DATA = 12'b000000000100;
            14'b00_101111011010: DATA = 12'b000000000100;
            14'b00_101111011011: DATA = 12'b000000000100;
            14'b00_101111011100: DATA = 12'b000000000100;
            14'b00_101111011101: DATA = 12'b000000000011;
            14'b00_101111011110: DATA = 12'b000000000011;
            14'b00_101111011111: DATA = 12'b000000000011;
            14'b00_101111100000: DATA = 12'b000000000011;
            14'b00_101111100001: DATA = 12'b000000000011;
            14'b00_101111100010: DATA = 12'b000000000011;
            14'b00_101111100011: DATA = 12'b000000000011;
            14'b00_101111100100: DATA = 12'b000000000010;
            14'b00_101111100101: DATA = 12'b000000000010;
            14'b00_101111100110: DATA = 12'b000000000010;
            14'b00_101111100111: DATA = 12'b000000000010;
            14'b00_101111101000: DATA = 12'b000000000010;
            14'b00_101111101001: DATA = 12'b000000000010;
            14'b00_101111101010: DATA = 12'b000000000010;
            14'b00_101111101011: DATA = 12'b000000000010;
            14'b00_101111101100: DATA = 12'b000000000001;
            14'b00_101111101101: DATA = 12'b000000000001;
            14'b00_101111101110: DATA = 12'b000000000001;
            14'b00_101111101111: DATA = 12'b000000000001;
            14'b00_101111110000: DATA = 12'b000000000001;
            14'b00_101111110001: DATA = 12'b000000000001;
            14'b00_101111110010: DATA = 12'b000000000001;
            14'b00_101111110011: DATA = 12'b000000000001;
            14'b00_101111110100: DATA = 12'b000000000001;
            14'b00_101111110101: DATA = 12'b000000000001;
            14'b00_101111110110: DATA = 12'b000000000001;
            14'b00_101111110111: DATA = 12'b000000000001;
            14'b00_101111111000: DATA = 12'b000000000001;
            14'b00_101111111001: DATA = 12'b000000000001;
            14'b00_101111111010: DATA = 12'b000000000001;
            14'b00_101111111011: DATA = 12'b000000000001;
            14'b00_101111111100: DATA = 12'b000000000001;
            14'b00_101111111101: DATA = 12'b000000000001;
            14'b00_101111111110: DATA = 12'b000000000001;
            14'b00_101111111111: DATA = 12'b000000000001;
            14'b00_110000000000: DATA = 12'b000000000001;
            14'b00_110000000001: DATA = 12'b000000000001;
            14'b00_110000000010: DATA = 12'b000000000001;
            14'b00_110000000011: DATA = 12'b000000000001;
            14'b00_110000000100: DATA = 12'b000000000001;
            14'b00_110000000101: DATA = 12'b000000000001;
            14'b00_110000000110: DATA = 12'b000000000001;
            14'b00_110000000111: DATA = 12'b000000000001;
            14'b00_110000001000: DATA = 12'b000000000001;
            14'b00_110000001001: DATA = 12'b000000000001;
            14'b00_110000001010: DATA = 12'b000000000001;
            14'b00_110000001011: DATA = 12'b000000000001;
            14'b00_110000001100: DATA = 12'b000000000001;
            14'b00_110000001101: DATA = 12'b000000000001;
            14'b00_110000001110: DATA = 12'b000000000001;
            14'b00_110000001111: DATA = 12'b000000000001;
            14'b00_110000010000: DATA = 12'b000000000001;
            14'b00_110000010001: DATA = 12'b000000000001;
            14'b00_110000010010: DATA = 12'b000000000001;
            14'b00_110000010011: DATA = 12'b000000000001;
            14'b00_110000010100: DATA = 12'b000000000001;
            14'b00_110000010101: DATA = 12'b000000000010;
            14'b00_110000010110: DATA = 12'b000000000010;
            14'b00_110000010111: DATA = 12'b000000000010;
            14'b00_110000011000: DATA = 12'b000000000010;
            14'b00_110000011001: DATA = 12'b000000000010;
            14'b00_110000011010: DATA = 12'b000000000010;
            14'b00_110000011011: DATA = 12'b000000000010;
            14'b00_110000011100: DATA = 12'b000000000010;
            14'b00_110000011101: DATA = 12'b000000000011;
            14'b00_110000011110: DATA = 12'b000000000011;
            14'b00_110000011111: DATA = 12'b000000000011;
            14'b00_110000100000: DATA = 12'b000000000011;
            14'b00_110000100001: DATA = 12'b000000000011;
            14'b00_110000100010: DATA = 12'b000000000011;
            14'b00_110000100011: DATA = 12'b000000000011;
            14'b00_110000100100: DATA = 12'b000000000100;
            14'b00_110000100101: DATA = 12'b000000000100;
            14'b00_110000100110: DATA = 12'b000000000100;
            14'b00_110000100111: DATA = 12'b000000000100;
            14'b00_110000101000: DATA = 12'b000000000100;
            14'b00_110000101001: DATA = 12'b000000000101;
            14'b00_110000101010: DATA = 12'b000000000101;
            14'b00_110000101011: DATA = 12'b000000000101;
            14'b00_110000101100: DATA = 12'b000000000101;
            14'b00_110000101101: DATA = 12'b000000000101;
            14'b00_110000101110: DATA = 12'b000000000110;
            14'b00_110000101111: DATA = 12'b000000000110;
            14'b00_110000110000: DATA = 12'b000000000110;
            14'b00_110000110001: DATA = 12'b000000000110;
            14'b00_110000110010: DATA = 12'b000000000111;
            14'b00_110000110011: DATA = 12'b000000000111;
            14'b00_110000110100: DATA = 12'b000000000111;
            14'b00_110000110101: DATA = 12'b000000000111;
            14'b00_110000110110: DATA = 12'b000000001000;
            14'b00_110000110111: DATA = 12'b000000001000;
            14'b00_110000111000: DATA = 12'b000000001000;
            14'b00_110000111001: DATA = 12'b000000001000;
            14'b00_110000111010: DATA = 12'b000000001001;
            14'b00_110000111011: DATA = 12'b000000001001;
            14'b00_110000111100: DATA = 12'b000000001001;
            14'b00_110000111101: DATA = 12'b000000001001;
            14'b00_110000111110: DATA = 12'b000000001010;
            14'b00_110000111111: DATA = 12'b000000001010;
            14'b00_110001000000: DATA = 12'b000000001010;
            14'b00_110001000001: DATA = 12'b000000001011;
            14'b00_110001000010: DATA = 12'b000000001011;
            14'b00_110001000011: DATA = 12'b000000001011;
            14'b00_110001000100: DATA = 12'b000000001100;
            14'b00_110001000101: DATA = 12'b000000001100;
            14'b00_110001000110: DATA = 12'b000000001100;
            14'b00_110001000111: DATA = 12'b000000001101;
            14'b00_110001001000: DATA = 12'b000000001101;
            14'b00_110001001001: DATA = 12'b000000001101;
            14'b00_110001001010: DATA = 12'b000000001110;
            14'b00_110001001011: DATA = 12'b000000001110;
            14'b00_110001001100: DATA = 12'b000000001110;
            14'b00_110001001101: DATA = 12'b000000001111;
            14'b00_110001001110: DATA = 12'b000000001111;
            14'b00_110001001111: DATA = 12'b000000010000;
            14'b00_110001010000: DATA = 12'b000000010000;
            14'b00_110001010001: DATA = 12'b000000010000;
            14'b00_110001010010: DATA = 12'b000000010001;
            14'b00_110001010011: DATA = 12'b000000010001;
            14'b00_110001010100: DATA = 12'b000000010001;
            14'b00_110001010101: DATA = 12'b000000010010;
            14'b00_110001010110: DATA = 12'b000000010010;
            14'b00_110001010111: DATA = 12'b000000010011;
            14'b00_110001011000: DATA = 12'b000000010011;
            14'b00_110001011001: DATA = 12'b000000010100;
            14'b00_110001011010: DATA = 12'b000000010100;
            14'b00_110001011011: DATA = 12'b000000010100;
            14'b00_110001011100: DATA = 12'b000000010101;
            14'b00_110001011101: DATA = 12'b000000010101;
            14'b00_110001011110: DATA = 12'b000000010110;
            14'b00_110001011111: DATA = 12'b000000010110;
            14'b00_110001100000: DATA = 12'b000000010111;
            14'b00_110001100001: DATA = 12'b000000010111;
            14'b00_110001100010: DATA = 12'b000000011000;
            14'b00_110001100011: DATA = 12'b000000011000;
            14'b00_110001100100: DATA = 12'b000000011001;
            14'b00_110001100101: DATA = 12'b000000011001;
            14'b00_110001100110: DATA = 12'b000000011010;
            14'b00_110001100111: DATA = 12'b000000011010;
            14'b00_110001101000: DATA = 12'b000000011010;
            14'b00_110001101001: DATA = 12'b000000011011;
            14'b00_110001101010: DATA = 12'b000000011100;
            14'b00_110001101011: DATA = 12'b000000011100;
            14'b00_110001101100: DATA = 12'b000000011101;
            14'b00_110001101101: DATA = 12'b000000011101;
            14'b00_110001101110: DATA = 12'b000000011110;
            14'b00_110001101111: DATA = 12'b000000011110;
            14'b00_110001110000: DATA = 12'b000000011111;
            14'b00_110001110001: DATA = 12'b000000011111;
            14'b00_110001110010: DATA = 12'b000000100000;
            14'b00_110001110011: DATA = 12'b000000100000;
            14'b00_110001110100: DATA = 12'b000000100001;
            14'b00_110001110101: DATA = 12'b000000100001;
            14'b00_110001110110: DATA = 12'b000000100010;
            14'b00_110001110111: DATA = 12'b000000100011;
            14'b00_110001111000: DATA = 12'b000000100011;
            14'b00_110001111001: DATA = 12'b000000100100;
            14'b00_110001111010: DATA = 12'b000000100100;
            14'b00_110001111011: DATA = 12'b000000100101;
            14'b00_110001111100: DATA = 12'b000000100101;
            14'b00_110001111101: DATA = 12'b000000100110;
            14'b00_110001111110: DATA = 12'b000000100111;
            14'b00_110001111111: DATA = 12'b000000100111;
            14'b00_110010000000: DATA = 12'b000000101000;
            14'b00_110010000001: DATA = 12'b000000101000;
            14'b00_110010000010: DATA = 12'b000000101001;
            14'b00_110010000011: DATA = 12'b000000101010;
            14'b00_110010000100: DATA = 12'b000000101010;
            14'b00_110010000101: DATA = 12'b000000101011;
            14'b00_110010000110: DATA = 12'b000000101100;
            14'b00_110010000111: DATA = 12'b000000101100;
            14'b00_110010001000: DATA = 12'b000000101101;
            14'b00_110010001001: DATA = 12'b000000101110;
            14'b00_110010001010: DATA = 12'b000000101110;
            14'b00_110010001011: DATA = 12'b000000101111;
            14'b00_110010001100: DATA = 12'b000000110000;
            14'b00_110010001101: DATA = 12'b000000110000;
            14'b00_110010001110: DATA = 12'b000000110001;
            14'b00_110010001111: DATA = 12'b000000110010;
            14'b00_110010010000: DATA = 12'b000000110010;
            14'b00_110010010001: DATA = 12'b000000110011;
            14'b00_110010010010: DATA = 12'b000000110100;
            14'b00_110010010011: DATA = 12'b000000110100;
            14'b00_110010010100: DATA = 12'b000000110101;
            14'b00_110010010101: DATA = 12'b000000110110;
            14'b00_110010010110: DATA = 12'b000000110110;
            14'b00_110010010111: DATA = 12'b000000110111;
            14'b00_110010011000: DATA = 12'b000000111000;
            14'b00_110010011001: DATA = 12'b000000111001;
            14'b00_110010011010: DATA = 12'b000000111001;
            14'b00_110010011011: DATA = 12'b000000111010;
            14'b00_110010011100: DATA = 12'b000000111011;
            14'b00_110010011101: DATA = 12'b000000111100;
            14'b00_110010011110: DATA = 12'b000000111100;
            14'b00_110010011111: DATA = 12'b000000111101;
            14'b00_110010100000: DATA = 12'b000000111110;
            14'b00_110010100001: DATA = 12'b000000111111;
            14'b00_110010100010: DATA = 12'b000000111111;
            14'b00_110010100011: DATA = 12'b000001000000;
            14'b00_110010100100: DATA = 12'b000001000001;
            14'b00_110010100101: DATA = 12'b000001000010;
            14'b00_110010100110: DATA = 12'b000001000011;
            14'b00_110010100111: DATA = 12'b000001000011;
            14'b00_110010101000: DATA = 12'b000001000100;
            14'b00_110010101001: DATA = 12'b000001000101;
            14'b00_110010101010: DATA = 12'b000001000110;
            14'b00_110010101011: DATA = 12'b000001000111;
            14'b00_110010101100: DATA = 12'b000001000111;
            14'b00_110010101101: DATA = 12'b000001001000;
            14'b00_110010101110: DATA = 12'b000001001001;
            14'b00_110010101111: DATA = 12'b000001001010;
            14'b00_110010110000: DATA = 12'b000001001011;
            14'b00_110010110001: DATA = 12'b000001001011;
            14'b00_110010110010: DATA = 12'b000001001100;
            14'b00_110010110011: DATA = 12'b000001001101;
            14'b00_110010110100: DATA = 12'b000001001110;
            14'b00_110010110101: DATA = 12'b000001001111;
            14'b00_110010110110: DATA = 12'b000001010000;
            14'b00_110010110111: DATA = 12'b000001010001;
            14'b00_110010111000: DATA = 12'b000001010001;
            14'b00_110010111001: DATA = 12'b000001010010;
            14'b00_110010111010: DATA = 12'b000001010011;
            14'b00_110010111011: DATA = 12'b000001010100;
            14'b00_110010111100: DATA = 12'b000001010101;
            14'b00_110010111101: DATA = 12'b000001010110;
            14'b00_110010111110: DATA = 12'b000001010111;
            14'b00_110010111111: DATA = 12'b000001011000;
            14'b00_110011000000: DATA = 12'b000001011001;
            14'b00_110011000001: DATA = 12'b000001011010;
            14'b00_110011000010: DATA = 12'b000001011010;
            14'b00_110011000011: DATA = 12'b000001011011;
            14'b00_110011000100: DATA = 12'b000001011100;
            14'b00_110011000101: DATA = 12'b000001011101;
            14'b00_110011000110: DATA = 12'b000001011110;
            14'b00_110011000111: DATA = 12'b000001011111;
            14'b00_110011001000: DATA = 12'b000001100000;
            14'b00_110011001001: DATA = 12'b000001100001;
            14'b00_110011001010: DATA = 12'b000001100010;
            14'b00_110011001011: DATA = 12'b000001100011;
            14'b00_110011001100: DATA = 12'b000001100100;
            14'b00_110011001101: DATA = 12'b000001100101;
            14'b00_110011001110: DATA = 12'b000001100110;
            14'b00_110011001111: DATA = 12'b000001100111;
            14'b00_110011010000: DATA = 12'b000001101000;
            14'b00_110011010001: DATA = 12'b000001101001;
            14'b00_110011010010: DATA = 12'b000001101010;
            14'b00_110011010011: DATA = 12'b000001101011;
            14'b00_110011010100: DATA = 12'b000001101100;
            14'b00_110011010101: DATA = 12'b000001101101;
            14'b00_110011010110: DATA = 12'b000001101110;
            14'b00_110011010111: DATA = 12'b000001101111;
            14'b00_110011011000: DATA = 12'b000001110000;
            14'b00_110011011001: DATA = 12'b000001110001;
            14'b00_110011011010: DATA = 12'b000001110010;
            14'b00_110011011011: DATA = 12'b000001110011;
            14'b00_110011011100: DATA = 12'b000001110100;
            14'b00_110011011101: DATA = 12'b000001110101;
            14'b00_110011011110: DATA = 12'b000001110110;
            14'b00_110011011111: DATA = 12'b000001110111;
            14'b00_110011100000: DATA = 12'b000001111000;
            14'b00_110011100001: DATA = 12'b000001111001;
            14'b00_110011100010: DATA = 12'b000001111010;
            14'b00_110011100011: DATA = 12'b000001111011;
            14'b00_110011100100: DATA = 12'b000001111100;
            14'b00_110011100101: DATA = 12'b000001111110;
            14'b00_110011100110: DATA = 12'b000001111111;
            14'b00_110011100111: DATA = 12'b000010000000;
            14'b00_110011101000: DATA = 12'b000010000001;
            14'b00_110011101001: DATA = 12'b000010000010;
            14'b00_110011101010: DATA = 12'b000010000011;
            14'b00_110011101011: DATA = 12'b000010000100;
            14'b00_110011101100: DATA = 12'b000010000101;
            14'b00_110011101101: DATA = 12'b000010000110;
            14'b00_110011101110: DATA = 12'b000010000111;
            14'b00_110011101111: DATA = 12'b000010001001;
            14'b00_110011110000: DATA = 12'b000010001010;
            14'b00_110011110001: DATA = 12'b000010001011;
            14'b00_110011110010: DATA = 12'b000010001100;
            14'b00_110011110011: DATA = 12'b000010001101;
            14'b00_110011110100: DATA = 12'b000010001110;
            14'b00_110011110101: DATA = 12'b000010001111;
            14'b00_110011110110: DATA = 12'b000010010001;
            14'b00_110011110111: DATA = 12'b000010010010;
            14'b00_110011111000: DATA = 12'b000010010011;
            14'b00_110011111001: DATA = 12'b000010010100;
            14'b00_110011111010: DATA = 12'b000010010101;
            14'b00_110011111011: DATA = 12'b000010010110;
            14'b00_110011111100: DATA = 12'b000010011000;
            14'b00_110011111101: DATA = 12'b000010011001;
            14'b00_110011111110: DATA = 12'b000010011010;
            14'b00_110011111111: DATA = 12'b000010011011;
            14'b00_110100000000: DATA = 12'b000010011100;
            14'b00_110100000001: DATA = 12'b000010011110;
            14'b00_110100000010: DATA = 12'b000010011111;
            14'b00_110100000011: DATA = 12'b000010100000;
            14'b00_110100000100: DATA = 12'b000010100001;
            14'b00_110100000101: DATA = 12'b000010100010;
            14'b00_110100000110: DATA = 12'b000010100100;
            14'b00_110100000111: DATA = 12'b000010100101;
            14'b00_110100001000: DATA = 12'b000010100110;
            14'b00_110100001001: DATA = 12'b000010100111;
            14'b00_110100001010: DATA = 12'b000010101001;
            14'b00_110100001011: DATA = 12'b000010101010;
            14'b00_110100001100: DATA = 12'b000010101011;
            14'b00_110100001101: DATA = 12'b000010101100;
            14'b00_110100001110: DATA = 12'b000010101110;
            14'b00_110100001111: DATA = 12'b000010101111;
            14'b00_110100010000: DATA = 12'b000010110000;
            14'b00_110100010001: DATA = 12'b000010110001;
            14'b00_110100010010: DATA = 12'b000010110011;
            14'b00_110100010011: DATA = 12'b000010110100;
            14'b00_110100010100: DATA = 12'b000010110101;
            14'b00_110100010101: DATA = 12'b000010110111;
            14'b00_110100010110: DATA = 12'b000010111000;
            14'b00_110100010111: DATA = 12'b000010111001;
            14'b00_110100011000: DATA = 12'b000010111010;
            14'b00_110100011001: DATA = 12'b000010111100;
            14'b00_110100011010: DATA = 12'b000010111101;
            14'b00_110100011011: DATA = 12'b000010111110;
            14'b00_110100011100: DATA = 12'b000011000000;
            14'b00_110100011101: DATA = 12'b000011000001;
            14'b00_110100011110: DATA = 12'b000011000010;
            14'b00_110100011111: DATA = 12'b000011000100;
            14'b00_110100100000: DATA = 12'b000011000101;
            14'b00_110100100001: DATA = 12'b000011000110;
            14'b00_110100100010: DATA = 12'b000011001000;
            14'b00_110100100011: DATA = 12'b000011001001;
            14'b00_110100100100: DATA = 12'b000011001010;
            14'b00_110100100101: DATA = 12'b000011001100;
            14'b00_110100100110: DATA = 12'b000011001101;
            14'b00_110100100111: DATA = 12'b000011001111;
            14'b00_110100101000: DATA = 12'b000011010000;
            14'b00_110100101001: DATA = 12'b000011010001;
            14'b00_110100101010: DATA = 12'b000011010011;
            14'b00_110100101011: DATA = 12'b000011010100;
            14'b00_110100101100: DATA = 12'b000011010101;
            14'b00_110100101101: DATA = 12'b000011010111;
            14'b00_110100101110: DATA = 12'b000011011000;
            14'b00_110100101111: DATA = 12'b000011011010;
            14'b00_110100110000: DATA = 12'b000011011011;
            14'b00_110100110001: DATA = 12'b000011011100;
            14'b00_110100110010: DATA = 12'b000011011110;
            14'b00_110100110011: DATA = 12'b000011011111;
            14'b00_110100110100: DATA = 12'b000011100001;
            14'b00_110100110101: DATA = 12'b000011100010;
            14'b00_110100110110: DATA = 12'b000011100100;
            14'b00_110100110111: DATA = 12'b000011100101;
            14'b00_110100111000: DATA = 12'b000011100111;
            14'b00_110100111001: DATA = 12'b000011101000;
            14'b00_110100111010: DATA = 12'b000011101001;
            14'b00_110100111011: DATA = 12'b000011101011;
            14'b00_110100111100: DATA = 12'b000011101100;
            14'b00_110100111101: DATA = 12'b000011101110;
            14'b00_110100111110: DATA = 12'b000011101111;
            14'b00_110100111111: DATA = 12'b000011110001;
            14'b00_110101000000: DATA = 12'b000011110010;
            14'b00_110101000001: DATA = 12'b000011110100;
            14'b00_110101000010: DATA = 12'b000011110101;
            14'b00_110101000011: DATA = 12'b000011110111;
            14'b00_110101000100: DATA = 12'b000011111000;
            14'b00_110101000101: DATA = 12'b000011111010;
            14'b00_110101000110: DATA = 12'b000011111011;
            14'b00_110101000111: DATA = 12'b000011111101;
            14'b00_110101001000: DATA = 12'b000011111110;
            14'b00_110101001001: DATA = 12'b000100000000;
            14'b00_110101001010: DATA = 12'b000100000001;
            14'b00_110101001011: DATA = 12'b000100000011;
            14'b00_110101001100: DATA = 12'b000100000100;
            14'b00_110101001101: DATA = 12'b000100000110;
            14'b00_110101001110: DATA = 12'b000100000111;
            14'b00_110101001111: DATA = 12'b000100001001;
            14'b00_110101010000: DATA = 12'b000100001010;
            14'b00_110101010001: DATA = 12'b000100001100;
            14'b00_110101010010: DATA = 12'b000100001110;
            14'b00_110101010011: DATA = 12'b000100001111;
            14'b00_110101010100: DATA = 12'b000100010001;
            14'b00_110101010101: DATA = 12'b000100010010;
            14'b00_110101010110: DATA = 12'b000100010100;
            14'b00_110101010111: DATA = 12'b000100010101;
            14'b00_110101011000: DATA = 12'b000100010111;
            14'b00_110101011001: DATA = 12'b000100011001;
            14'b00_110101011010: DATA = 12'b000100011010;
            14'b00_110101011011: DATA = 12'b000100011100;
            14'b00_110101011100: DATA = 12'b000100011101;
            14'b00_110101011101: DATA = 12'b000100011111;
            14'b00_110101011110: DATA = 12'b000100100001;
            14'b00_110101011111: DATA = 12'b000100100010;
            14'b00_110101100000: DATA = 12'b000100100100;
            14'b00_110101100001: DATA = 12'b000100100101;
            14'b00_110101100010: DATA = 12'b000100100111;
            14'b00_110101100011: DATA = 12'b000100101001;
            14'b00_110101100100: DATA = 12'b000100101010;
            14'b00_110101100101: DATA = 12'b000100101100;
            14'b00_110101100110: DATA = 12'b000100101101;
            14'b00_110101100111: DATA = 12'b000100101111;
            14'b00_110101101000: DATA = 12'b000100110001;
            14'b00_110101101001: DATA = 12'b000100110010;
            14'b00_110101101010: DATA = 12'b000100110100;
            14'b00_110101101011: DATA = 12'b000100110110;
            14'b00_110101101100: DATA = 12'b000100110111;
            14'b00_110101101101: DATA = 12'b000100111001;
            14'b00_110101101110: DATA = 12'b000100111011;
            14'b00_110101101111: DATA = 12'b000100111100;
            14'b00_110101110000: DATA = 12'b000100111110;
            14'b00_110101110001: DATA = 12'b000101000000;
            14'b00_110101110010: DATA = 12'b000101000001;
            14'b00_110101110011: DATA = 12'b000101000011;
            14'b00_110101110100: DATA = 12'b000101000101;
            14'b00_110101110101: DATA = 12'b000101000111;
            14'b00_110101110110: DATA = 12'b000101001000;
            14'b00_110101110111: DATA = 12'b000101001010;
            14'b00_110101111000: DATA = 12'b000101001100;
            14'b00_110101111001: DATA = 12'b000101001101;
            14'b00_110101111010: DATA = 12'b000101001111;
            14'b00_110101111011: DATA = 12'b000101010001;
            14'b00_110101111100: DATA = 12'b000101010011;
            14'b00_110101111101: DATA = 12'b000101010100;
            14'b00_110101111110: DATA = 12'b000101010110;
            14'b00_110101111111: DATA = 12'b000101011000;
            14'b00_110110000000: DATA = 12'b000101011001;
            14'b00_110110000001: DATA = 12'b000101011011;
            14'b00_110110000010: DATA = 12'b000101011101;
            14'b00_110110000011: DATA = 12'b000101011111;
            14'b00_110110000100: DATA = 12'b000101100000;
            14'b00_110110000101: DATA = 12'b000101100010;
            14'b00_110110000110: DATA = 12'b000101100100;
            14'b00_110110000111: DATA = 12'b000101100110;
            14'b00_110110001000: DATA = 12'b000101101000;
            14'b00_110110001001: DATA = 12'b000101101001;
            14'b00_110110001010: DATA = 12'b000101101011;
            14'b00_110110001011: DATA = 12'b000101101101;
            14'b00_110110001100: DATA = 12'b000101101111;
            14'b00_110110001101: DATA = 12'b000101110000;
            14'b00_110110001110: DATA = 12'b000101110010;
            14'b00_110110001111: DATA = 12'b000101110100;
            14'b00_110110010000: DATA = 12'b000101110110;
            14'b00_110110010001: DATA = 12'b000101111000;
            14'b00_110110010010: DATA = 12'b000101111010;
            14'b00_110110010011: DATA = 12'b000101111011;
            14'b00_110110010100: DATA = 12'b000101111101;
            14'b00_110110010101: DATA = 12'b000101111111;
            14'b00_110110010110: DATA = 12'b000110000001;
            14'b00_110110010111: DATA = 12'b000110000011;
            14'b00_110110011000: DATA = 12'b000110000100;
            14'b00_110110011001: DATA = 12'b000110000110;
            14'b00_110110011010: DATA = 12'b000110001000;
            14'b00_110110011011: DATA = 12'b000110001010;
            14'b00_110110011100: DATA = 12'b000110001100;
            14'b00_110110011101: DATA = 12'b000110001110;
            14'b00_110110011110: DATA = 12'b000110010000;
            14'b00_110110011111: DATA = 12'b000110010001;
            14'b00_110110100000: DATA = 12'b000110010011;
            14'b00_110110100001: DATA = 12'b000110010101;
            14'b00_110110100010: DATA = 12'b000110010111;
            14'b00_110110100011: DATA = 12'b000110011001;
            14'b00_110110100100: DATA = 12'b000110011011;
            14'b00_110110100101: DATA = 12'b000110011101;
            14'b00_110110100110: DATA = 12'b000110011111;
            14'b00_110110100111: DATA = 12'b000110100001;
            14'b00_110110101000: DATA = 12'b000110100010;
            14'b00_110110101001: DATA = 12'b000110100100;
            14'b00_110110101010: DATA = 12'b000110100110;
            14'b00_110110101011: DATA = 12'b000110101000;
            14'b00_110110101100: DATA = 12'b000110101010;
            14'b00_110110101101: DATA = 12'b000110101100;
            14'b00_110110101110: DATA = 12'b000110101110;
            14'b00_110110101111: DATA = 12'b000110110000;
            14'b00_110110110000: DATA = 12'b000110110010;
            14'b00_110110110001: DATA = 12'b000110110100;
            14'b00_110110110010: DATA = 12'b000110110110;
            14'b00_110110110011: DATA = 12'b000110111000;
            14'b00_110110110100: DATA = 12'b000110111010;
            14'b00_110110110101: DATA = 12'b000110111011;
            14'b00_110110110110: DATA = 12'b000110111101;
            14'b00_110110110111: DATA = 12'b000110111111;
            14'b00_110110111000: DATA = 12'b000111000001;
            14'b00_110110111001: DATA = 12'b000111000011;
            14'b00_110110111010: DATA = 12'b000111000101;
            14'b00_110110111011: DATA = 12'b000111000111;
            14'b00_110110111100: DATA = 12'b000111001001;
            14'b00_110110111101: DATA = 12'b000111001011;
            14'b00_110110111110: DATA = 12'b000111001101;
            14'b00_110110111111: DATA = 12'b000111001111;
            14'b00_110111000000: DATA = 12'b000111010001;
            14'b00_110111000001: DATA = 12'b000111010011;
            14'b00_110111000010: DATA = 12'b000111010101;
            14'b00_110111000011: DATA = 12'b000111010111;
            14'b00_110111000100: DATA = 12'b000111011001;
            14'b00_110111000101: DATA = 12'b000111011011;
            14'b00_110111000110: DATA = 12'b000111011101;
            14'b00_110111000111: DATA = 12'b000111011111;
            14'b00_110111001000: DATA = 12'b000111100001;
            14'b00_110111001001: DATA = 12'b000111100011;
            14'b00_110111001010: DATA = 12'b000111100101;
            14'b00_110111001011: DATA = 12'b000111100111;
            14'b00_110111001100: DATA = 12'b000111101001;
            14'b00_110111001101: DATA = 12'b000111101011;
            14'b00_110111001110: DATA = 12'b000111101101;
            14'b00_110111001111: DATA = 12'b000111101111;
            14'b00_110111010000: DATA = 12'b000111110001;
            14'b00_110111010001: DATA = 12'b000111110100;
            14'b00_110111010010: DATA = 12'b000111110110;
            14'b00_110111010011: DATA = 12'b000111111000;
            14'b00_110111010100: DATA = 12'b000111111010;
            14'b00_110111010101: DATA = 12'b000111111100;
            14'b00_110111010110: DATA = 12'b000111111110;
            14'b00_110111010111: DATA = 12'b001000000000;
            14'b00_110111011000: DATA = 12'b001000000010;
            14'b00_110111011001: DATA = 12'b001000000100;
            14'b00_110111011010: DATA = 12'b001000000110;
            14'b00_110111011011: DATA = 12'b001000001000;
            14'b00_110111011100: DATA = 12'b001000001010;
            14'b00_110111011101: DATA = 12'b001000001100;
            14'b00_110111011110: DATA = 12'b001000001111;
            14'b00_110111011111: DATA = 12'b001000010001;
            14'b00_110111100000: DATA = 12'b001000010011;
            14'b00_110111100001: DATA = 12'b001000010101;
            14'b00_110111100010: DATA = 12'b001000010111;
            14'b00_110111100011: DATA = 12'b001000011001;
            14'b00_110111100100: DATA = 12'b001000011011;
            14'b00_110111100101: DATA = 12'b001000011101;
            14'b00_110111100110: DATA = 12'b001000011111;
            14'b00_110111100111: DATA = 12'b001000100010;
            14'b00_110111101000: DATA = 12'b001000100100;
            14'b00_110111101001: DATA = 12'b001000100110;
            14'b00_110111101010: DATA = 12'b001000101000;
            14'b00_110111101011: DATA = 12'b001000101010;
            14'b00_110111101100: DATA = 12'b001000101100;
            14'b00_110111101101: DATA = 12'b001000101110;
            14'b00_110111101110: DATA = 12'b001000110001;
            14'b00_110111101111: DATA = 12'b001000110011;
            14'b00_110111110000: DATA = 12'b001000110101;
            14'b00_110111110001: DATA = 12'b001000110111;
            14'b00_110111110010: DATA = 12'b001000111001;
            14'b00_110111110011: DATA = 12'b001000111011;
            14'b00_110111110100: DATA = 12'b001000111110;
            14'b00_110111110101: DATA = 12'b001001000000;
            14'b00_110111110110: DATA = 12'b001001000010;
            14'b00_110111110111: DATA = 12'b001001000100;
            14'b00_110111111000: DATA = 12'b001001000110;
            14'b00_110111111001: DATA = 12'b001001001001;
            14'b00_110111111010: DATA = 12'b001001001011;
            14'b00_110111111011: DATA = 12'b001001001101;
            14'b00_110111111100: DATA = 12'b001001001111;
            14'b00_110111111101: DATA = 12'b001001010001;
            14'b00_110111111110: DATA = 12'b001001010100;
            14'b00_110111111111: DATA = 12'b001001010110;
            14'b00_111000000000: DATA = 12'b001001011000;
            14'b00_111000000001: DATA = 12'b001001011010;
            14'b00_111000000010: DATA = 12'b001001011100;
            14'b00_111000000011: DATA = 12'b001001011111;
            14'b00_111000000100: DATA = 12'b001001100001;
            14'b00_111000000101: DATA = 12'b001001100011;
            14'b00_111000000110: DATA = 12'b001001100101;
            14'b00_111000000111: DATA = 12'b001001101000;
            14'b00_111000001000: DATA = 12'b001001101010;
            14'b00_111000001001: DATA = 12'b001001101100;
            14'b00_111000001010: DATA = 12'b001001101110;
            14'b00_111000001011: DATA = 12'b001001110001;
            14'b00_111000001100: DATA = 12'b001001110011;
            14'b00_111000001101: DATA = 12'b001001110101;
            14'b00_111000001110: DATA = 12'b001001110111;
            14'b00_111000001111: DATA = 12'b001001111010;
            14'b00_111000010000: DATA = 12'b001001111100;
            14'b00_111000010001: DATA = 12'b001001111110;
            14'b00_111000010010: DATA = 12'b001010000001;
            14'b00_111000010011: DATA = 12'b001010000011;
            14'b00_111000010100: DATA = 12'b001010000101;
            14'b00_111000010101: DATA = 12'b001010000111;
            14'b00_111000010110: DATA = 12'b001010001010;
            14'b00_111000010111: DATA = 12'b001010001100;
            14'b00_111000011000: DATA = 12'b001010001110;
            14'b00_111000011001: DATA = 12'b001010010001;
            14'b00_111000011010: DATA = 12'b001010010011;
            14'b00_111000011011: DATA = 12'b001010010101;
            14'b00_111000011100: DATA = 12'b001010011000;
            14'b00_111000011101: DATA = 12'b001010011010;
            14'b00_111000011110: DATA = 12'b001010011100;
            14'b00_111000011111: DATA = 12'b001010011110;
            14'b00_111000100000: DATA = 12'b001010100001;
            14'b00_111000100001: DATA = 12'b001010100011;
            14'b00_111000100010: DATA = 12'b001010100101;
            14'b00_111000100011: DATA = 12'b001010101000;
            14'b00_111000100100: DATA = 12'b001010101010;
            14'b00_111000100101: DATA = 12'b001010101100;
            14'b00_111000100110: DATA = 12'b001010101111;
            14'b00_111000100111: DATA = 12'b001010110001;
            14'b00_111000101000: DATA = 12'b001010110100;
            14'b00_111000101001: DATA = 12'b001010110110;
            14'b00_111000101010: DATA = 12'b001010111000;
            14'b00_111000101011: DATA = 12'b001010111011;
            14'b00_111000101100: DATA = 12'b001010111101;
            14'b00_111000101101: DATA = 12'b001010111111;
            14'b00_111000101110: DATA = 12'b001011000010;
            14'b00_111000101111: DATA = 12'b001011000100;
            14'b00_111000110000: DATA = 12'b001011000110;
            14'b00_111000110001: DATA = 12'b001011001001;
            14'b00_111000110010: DATA = 12'b001011001011;
            14'b00_111000110011: DATA = 12'b001011001110;
            14'b00_111000110100: DATA = 12'b001011010000;
            14'b00_111000110101: DATA = 12'b001011010010;
            14'b00_111000110110: DATA = 12'b001011010101;
            14'b00_111000110111: DATA = 12'b001011010111;
            14'b00_111000111000: DATA = 12'b001011011010;
            14'b00_111000111001: DATA = 12'b001011011100;
            14'b00_111000111010: DATA = 12'b001011011110;
            14'b00_111000111011: DATA = 12'b001011100001;
            14'b00_111000111100: DATA = 12'b001011100011;
            14'b00_111000111101: DATA = 12'b001011100110;
            14'b00_111000111110: DATA = 12'b001011101000;
            14'b00_111000111111: DATA = 12'b001011101010;
            14'b00_111001000000: DATA = 12'b001011101101;
            14'b00_111001000001: DATA = 12'b001011101111;
            14'b00_111001000010: DATA = 12'b001011110010;
            14'b00_111001000011: DATA = 12'b001011110100;
            14'b00_111001000100: DATA = 12'b001011110111;
            14'b00_111001000101: DATA = 12'b001011111001;
            14'b00_111001000110: DATA = 12'b001011111100;
            14'b00_111001000111: DATA = 12'b001011111110;
            14'b00_111001001000: DATA = 12'b001100000000;
            14'b00_111001001001: DATA = 12'b001100000011;
            14'b00_111001001010: DATA = 12'b001100000101;
            14'b00_111001001011: DATA = 12'b001100001000;
            14'b00_111001001100: DATA = 12'b001100001010;
            14'b00_111001001101: DATA = 12'b001100001101;
            14'b00_111001001110: DATA = 12'b001100001111;
            14'b00_111001001111: DATA = 12'b001100010010;
            14'b00_111001010000: DATA = 12'b001100010100;
            14'b00_111001010001: DATA = 12'b001100010111;
            14'b00_111001010010: DATA = 12'b001100011001;
            14'b00_111001010011: DATA = 12'b001100011100;
            14'b00_111001010100: DATA = 12'b001100011110;
            14'b00_111001010101: DATA = 12'b001100100001;
            14'b00_111001010110: DATA = 12'b001100100011;
            14'b00_111001010111: DATA = 12'b001100100110;
            14'b00_111001011000: DATA = 12'b001100101000;
            14'b00_111001011001: DATA = 12'b001100101011;
            14'b00_111001011010: DATA = 12'b001100101101;
            14'b00_111001011011: DATA = 12'b001100110000;
            14'b00_111001011100: DATA = 12'b001100110010;
            14'b00_111001011101: DATA = 12'b001100110101;
            14'b00_111001011110: DATA = 12'b001100110111;
            14'b00_111001011111: DATA = 12'b001100111010;
            14'b00_111001100000: DATA = 12'b001100111100;
            14'b00_111001100001: DATA = 12'b001100111111;
            14'b00_111001100010: DATA = 12'b001101000001;
            14'b00_111001100011: DATA = 12'b001101000100;
            14'b00_111001100100: DATA = 12'b001101000110;
            14'b00_111001100101: DATA = 12'b001101001001;
            14'b00_111001100110: DATA = 12'b001101001011;
            14'b00_111001100111: DATA = 12'b001101001110;
            14'b00_111001101000: DATA = 12'b001101010000;
            14'b00_111001101001: DATA = 12'b001101010011;
            14'b00_111001101010: DATA = 12'b001101010101;
            14'b00_111001101011: DATA = 12'b001101011000;
            14'b00_111001101100: DATA = 12'b001101011011;
            14'b00_111001101101: DATA = 12'b001101011101;
            14'b00_111001101110: DATA = 12'b001101100000;
            14'b00_111001101111: DATA = 12'b001101100010;
            14'b00_111001110000: DATA = 12'b001101100101;
            14'b00_111001110001: DATA = 12'b001101100111;
            14'b00_111001110010: DATA = 12'b001101101010;
            14'b00_111001110011: DATA = 12'b001101101101;
            14'b00_111001110100: DATA = 12'b001101101111;
            14'b00_111001110101: DATA = 12'b001101110010;
            14'b00_111001110110: DATA = 12'b001101110100;
            14'b00_111001110111: DATA = 12'b001101110111;
            14'b00_111001111000: DATA = 12'b001101111001;
            14'b00_111001111001: DATA = 12'b001101111100;
            14'b00_111001111010: DATA = 12'b001101111111;
            14'b00_111001111011: DATA = 12'b001110000001;
            14'b00_111001111100: DATA = 12'b001110000100;
            14'b00_111001111101: DATA = 12'b001110000110;
            14'b00_111001111110: DATA = 12'b001110001001;
            14'b00_111001111111: DATA = 12'b001110001100;
            14'b00_111010000000: DATA = 12'b001110001110;
            14'b00_111010000001: DATA = 12'b001110010001;
            14'b00_111010000010: DATA = 12'b001110010011;
            14'b00_111010000011: DATA = 12'b001110010110;
            14'b00_111010000100: DATA = 12'b001110011001;
            14'b00_111010000101: DATA = 12'b001110011011;
            14'b00_111010000110: DATA = 12'b001110011110;
            14'b00_111010000111: DATA = 12'b001110100001;
            14'b00_111010001000: DATA = 12'b001110100011;
            14'b00_111010001001: DATA = 12'b001110100110;
            14'b00_111010001010: DATA = 12'b001110101000;
            14'b00_111010001011: DATA = 12'b001110101011;
            14'b00_111010001100: DATA = 12'b001110101110;
            14'b00_111010001101: DATA = 12'b001110110000;
            14'b00_111010001110: DATA = 12'b001110110011;
            14'b00_111010001111: DATA = 12'b001110110110;
            14'b00_111010010000: DATA = 12'b001110111000;
            14'b00_111010010001: DATA = 12'b001110111011;
            14'b00_111010010010: DATA = 12'b001110111110;
            14'b00_111010010011: DATA = 12'b001111000000;
            14'b00_111010010100: DATA = 12'b001111000011;
            14'b00_111010010101: DATA = 12'b001111000110;
            14'b00_111010010110: DATA = 12'b001111001000;
            14'b00_111010010111: DATA = 12'b001111001011;
            14'b00_111010011000: DATA = 12'b001111001110;
            14'b00_111010011001: DATA = 12'b001111010000;
            14'b00_111010011010: DATA = 12'b001111010011;
            14'b00_111010011011: DATA = 12'b001111010110;
            14'b00_111010011100: DATA = 12'b001111011000;
            14'b00_111010011101: DATA = 12'b001111011011;
            14'b00_111010011110: DATA = 12'b001111011110;
            14'b00_111010011111: DATA = 12'b001111100000;
            14'b00_111010100000: DATA = 12'b001111100011;
            14'b00_111010100001: DATA = 12'b001111100110;
            14'b00_111010100010: DATA = 12'b001111101001;
            14'b00_111010100011: DATA = 12'b001111101011;
            14'b00_111010100100: DATA = 12'b001111101110;
            14'b00_111010100101: DATA = 12'b001111110001;
            14'b00_111010100110: DATA = 12'b001111110011;
            14'b00_111010100111: DATA = 12'b001111110110;
            14'b00_111010101000: DATA = 12'b001111111001;
            14'b00_111010101001: DATA = 12'b001111111011;
            14'b00_111010101010: DATA = 12'b001111111110;
            14'b00_111010101011: DATA = 12'b010000000001;
            14'b00_111010101100: DATA = 12'b010000000100;
            14'b00_111010101101: DATA = 12'b010000000110;
            14'b00_111010101110: DATA = 12'b010000001001;
            14'b00_111010101111: DATA = 12'b010000001100;
            14'b00_111010110000: DATA = 12'b010000001111;
            14'b00_111010110001: DATA = 12'b010000010001;
            14'b00_111010110010: DATA = 12'b010000010100;
            14'b00_111010110011: DATA = 12'b010000010111;
            14'b00_111010110100: DATA = 12'b010000011001;
            14'b00_111010110101: DATA = 12'b010000011100;
            14'b00_111010110110: DATA = 12'b010000011111;
            14'b00_111010110111: DATA = 12'b010000100010;
            14'b00_111010111000: DATA = 12'b010000100100;
            14'b00_111010111001: DATA = 12'b010000100111;
            14'b00_111010111010: DATA = 12'b010000101010;
            14'b00_111010111011: DATA = 12'b010000101101;
            14'b00_111010111100: DATA = 12'b010000101111;
            14'b00_111010111101: DATA = 12'b010000110010;
            14'b00_111010111110: DATA = 12'b010000110101;
            14'b00_111010111111: DATA = 12'b010000111000;
            14'b00_111011000000: DATA = 12'b010000111011;
            14'b00_111011000001: DATA = 12'b010000111101;
            14'b00_111011000010: DATA = 12'b010001000000;
            14'b00_111011000011: DATA = 12'b010001000011;
            14'b00_111011000100: DATA = 12'b010001000110;
            14'b00_111011000101: DATA = 12'b010001001000;
            14'b00_111011000110: DATA = 12'b010001001011;
            14'b00_111011000111: DATA = 12'b010001001110;
            14'b00_111011001000: DATA = 12'b010001010001;
            14'b00_111011001001: DATA = 12'b010001010100;
            14'b00_111011001010: DATA = 12'b010001010110;
            14'b00_111011001011: DATA = 12'b010001011001;
            14'b00_111011001100: DATA = 12'b010001011100;
            14'b00_111011001101: DATA = 12'b010001011111;
            14'b00_111011001110: DATA = 12'b010001100010;
            14'b00_111011001111: DATA = 12'b010001100100;
            14'b00_111011010000: DATA = 12'b010001100111;
            14'b00_111011010001: DATA = 12'b010001101010;
            14'b00_111011010010: DATA = 12'b010001101101;
            14'b00_111011010011: DATA = 12'b010001110000;
            14'b00_111011010100: DATA = 12'b010001110010;
            14'b00_111011010101: DATA = 12'b010001110101;
            14'b00_111011010110: DATA = 12'b010001111000;
            14'b00_111011010111: DATA = 12'b010001111011;
            14'b00_111011011000: DATA = 12'b010001111110;
            14'b00_111011011001: DATA = 12'b010010000000;
            14'b00_111011011010: DATA = 12'b010010000011;
            14'b00_111011011011: DATA = 12'b010010000110;
            14'b00_111011011100: DATA = 12'b010010001001;
            14'b00_111011011101: DATA = 12'b010010001100;
            14'b00_111011011110: DATA = 12'b010010001111;
            14'b00_111011011111: DATA = 12'b010010010001;
            14'b00_111011100000: DATA = 12'b010010010100;
            14'b00_111011100001: DATA = 12'b010010010111;
            14'b00_111011100010: DATA = 12'b010010011010;
            14'b00_111011100011: DATA = 12'b010010011101;
            14'b00_111011100100: DATA = 12'b010010100000;
            14'b00_111011100101: DATA = 12'b010010100011;
            14'b00_111011100110: DATA = 12'b010010100101;
            14'b00_111011100111: DATA = 12'b010010101000;
            14'b00_111011101000: DATA = 12'b010010101011;
            14'b00_111011101001: DATA = 12'b010010101110;
            14'b00_111011101010: DATA = 12'b010010110001;
            14'b00_111011101011: DATA = 12'b010010110100;
            14'b00_111011101100: DATA = 12'b010010110111;
            14'b00_111011101101: DATA = 12'b010010111001;
            14'b00_111011101110: DATA = 12'b010010111100;
            14'b00_111011101111: DATA = 12'b010010111111;
            14'b00_111011110000: DATA = 12'b010011000010;
            14'b00_111011110001: DATA = 12'b010011000101;
            14'b00_111011110010: DATA = 12'b010011001000;
            14'b00_111011110011: DATA = 12'b010011001011;
            14'b00_111011110100: DATA = 12'b010011001101;
            14'b00_111011110101: DATA = 12'b010011010000;
            14'b00_111011110110: DATA = 12'b010011010011;
            14'b00_111011110111: DATA = 12'b010011010110;
            14'b00_111011111000: DATA = 12'b010011011001;
            14'b00_111011111001: DATA = 12'b010011011100;
            14'b00_111011111010: DATA = 12'b010011011111;
            14'b00_111011111011: DATA = 12'b010011100010;
            14'b00_111011111100: DATA = 12'b010011100101;
            14'b00_111011111101: DATA = 12'b010011100111;
            14'b00_111011111110: DATA = 12'b010011101010;
            14'b00_111011111111: DATA = 12'b010011101101;
            14'b00_111100000000: DATA = 12'b010011110000;
            14'b00_111100000001: DATA = 12'b010011110011;
            14'b00_111100000010: DATA = 12'b010011110110;
            14'b00_111100000011: DATA = 12'b010011111001;
            14'b00_111100000100: DATA = 12'b010011111100;
            14'b00_111100000101: DATA = 12'b010011111111;
            14'b00_111100000110: DATA = 12'b010100000010;
            14'b00_111100000111: DATA = 12'b010100000100;
            14'b00_111100001000: DATA = 12'b010100000111;
            14'b00_111100001001: DATA = 12'b010100001010;
            14'b00_111100001010: DATA = 12'b010100001101;
            14'b00_111100001011: DATA = 12'b010100010000;
            14'b00_111100001100: DATA = 12'b010100010011;
            14'b00_111100001101: DATA = 12'b010100010110;
            14'b00_111100001110: DATA = 12'b010100011001;
            14'b00_111100001111: DATA = 12'b010100011100;
            14'b00_111100010000: DATA = 12'b010100011111;
            14'b00_111100010001: DATA = 12'b010100100010;
            14'b00_111100010010: DATA = 12'b010100100101;
            14'b00_111100010011: DATA = 12'b010100101000;
            14'b00_111100010100: DATA = 12'b010100101011;
            14'b00_111100010101: DATA = 12'b010100101101;
            14'b00_111100010110: DATA = 12'b010100110000;
            14'b00_111100010111: DATA = 12'b010100110011;
            14'b00_111100011000: DATA = 12'b010100110110;
            14'b00_111100011001: DATA = 12'b010100111001;
            14'b00_111100011010: DATA = 12'b010100111100;
            14'b00_111100011011: DATA = 12'b010100111111;
            14'b00_111100011100: DATA = 12'b010101000010;
            14'b00_111100011101: DATA = 12'b010101000101;
            14'b00_111100011110: DATA = 12'b010101001000;
            14'b00_111100011111: DATA = 12'b010101001011;
            14'b00_111100100000: DATA = 12'b010101001110;
            14'b00_111100100001: DATA = 12'b010101010001;
            14'b00_111100100010: DATA = 12'b010101010100;
            14'b00_111100100011: DATA = 12'b010101010111;
            14'b00_111100100100: DATA = 12'b010101011010;
            14'b00_111100100101: DATA = 12'b010101011101;
            14'b00_111100100110: DATA = 12'b010101100000;
            14'b00_111100100111: DATA = 12'b010101100011;
            14'b00_111100101000: DATA = 12'b010101100110;
            14'b00_111100101001: DATA = 12'b010101101001;
            14'b00_111100101010: DATA = 12'b010101101100;
            14'b00_111100101011: DATA = 12'b010101101111;
            14'b00_111100101100: DATA = 12'b010101110001;
            14'b00_111100101101: DATA = 12'b010101110100;
            14'b00_111100101110: DATA = 12'b010101110111;
            14'b00_111100101111: DATA = 12'b010101111010;
            14'b00_111100110000: DATA = 12'b010101111101;
            14'b00_111100110001: DATA = 12'b010110000000;
            14'b00_111100110010: DATA = 12'b010110000011;
            14'b00_111100110011: DATA = 12'b010110000110;
            14'b00_111100110100: DATA = 12'b010110001001;
            14'b00_111100110101: DATA = 12'b010110001100;
            14'b00_111100110110: DATA = 12'b010110001111;
            14'b00_111100110111: DATA = 12'b010110010010;
            14'b00_111100111000: DATA = 12'b010110010101;
            14'b00_111100111001: DATA = 12'b010110011000;
            14'b00_111100111010: DATA = 12'b010110011011;
            14'b00_111100111011: DATA = 12'b010110011110;
            14'b00_111100111100: DATA = 12'b010110100001;
            14'b00_111100111101: DATA = 12'b010110100100;
            14'b00_111100111110: DATA = 12'b010110100111;
            14'b00_111100111111: DATA = 12'b010110101010;
            14'b00_111101000000: DATA = 12'b010110101101;
            14'b00_111101000001: DATA = 12'b010110110000;
            14'b00_111101000010: DATA = 12'b010110110011;
            14'b00_111101000011: DATA = 12'b010110110110;
            14'b00_111101000100: DATA = 12'b010110111001;
            14'b00_111101000101: DATA = 12'b010110111100;
            14'b00_111101000110: DATA = 12'b010110111111;
            14'b00_111101000111: DATA = 12'b010111000010;
            14'b00_111101001000: DATA = 12'b010111000101;
            14'b00_111101001001: DATA = 12'b010111001000;
            14'b00_111101001010: DATA = 12'b010111001011;
            14'b00_111101001011: DATA = 12'b010111001110;
            14'b00_111101001100: DATA = 12'b010111010001;
            14'b00_111101001101: DATA = 12'b010111010100;
            14'b00_111101001110: DATA = 12'b010111010111;
            14'b00_111101001111: DATA = 12'b010111011011;
            14'b00_111101010000: DATA = 12'b010111011110;
            14'b00_111101010001: DATA = 12'b010111100001;
            14'b00_111101010010: DATA = 12'b010111100100;
            14'b00_111101010011: DATA = 12'b010111100111;
            14'b00_111101010100: DATA = 12'b010111101010;
            14'b00_111101010101: DATA = 12'b010111101101;
            14'b00_111101010110: DATA = 12'b010111110000;
            14'b00_111101010111: DATA = 12'b010111110011;
            14'b00_111101011000: DATA = 12'b010111110110;
            14'b00_111101011001: DATA = 12'b010111111001;
            14'b00_111101011010: DATA = 12'b010111111100;
            14'b00_111101011011: DATA = 12'b010111111111;
            14'b00_111101011100: DATA = 12'b011000000010;
            14'b00_111101011101: DATA = 12'b011000000101;
            14'b00_111101011110: DATA = 12'b011000001000;
            14'b00_111101011111: DATA = 12'b011000001011;
            14'b00_111101100000: DATA = 12'b011000001110;
            14'b00_111101100001: DATA = 12'b011000010001;
            14'b00_111101100010: DATA = 12'b011000010100;
            14'b00_111101100011: DATA = 12'b011000010111;
            14'b00_111101100100: DATA = 12'b011000011010;
            14'b00_111101100101: DATA = 12'b011000011101;
            14'b00_111101100110: DATA = 12'b011000100000;
            14'b00_111101100111: DATA = 12'b011000100011;
            14'b00_111101101000: DATA = 12'b011000100111;
            14'b00_111101101001: DATA = 12'b011000101010;
            14'b00_111101101010: DATA = 12'b011000101101;
            14'b00_111101101011: DATA = 12'b011000110000;
            14'b00_111101101100: DATA = 12'b011000110011;
            14'b00_111101101101: DATA = 12'b011000110110;
            14'b00_111101101110: DATA = 12'b011000111001;
            14'b00_111101101111: DATA = 12'b011000111100;
            14'b00_111101110000: DATA = 12'b011000111111;
            14'b00_111101110001: DATA = 12'b011001000010;
            14'b00_111101110010: DATA = 12'b011001000101;
            14'b00_111101110011: DATA = 12'b011001001000;
            14'b00_111101110100: DATA = 12'b011001001011;
            14'b00_111101110101: DATA = 12'b011001001110;
            14'b00_111101110110: DATA = 12'b011001010001;
            14'b00_111101110111: DATA = 12'b011001010100;
            14'b00_111101111000: DATA = 12'b011001011000;
            14'b00_111101111001: DATA = 12'b011001011011;
            14'b00_111101111010: DATA = 12'b011001011110;
            14'b00_111101111011: DATA = 12'b011001100001;
            14'b00_111101111100: DATA = 12'b011001100100;
            14'b00_111101111101: DATA = 12'b011001100111;
            14'b00_111101111110: DATA = 12'b011001101010;
            14'b00_111101111111: DATA = 12'b011001101101;
            14'b00_111110000000: DATA = 12'b011001110000;
            14'b00_111110000001: DATA = 12'b011001110011;
            14'b00_111110000010: DATA = 12'b011001110110;
            14'b00_111110000011: DATA = 12'b011001111001;
            14'b00_111110000100: DATA = 12'b011001111100;
            14'b00_111110000101: DATA = 12'b011010000000;
            14'b00_111110000110: DATA = 12'b011010000011;
            14'b00_111110000111: DATA = 12'b011010000110;
            14'b00_111110001000: DATA = 12'b011010001001;
            14'b00_111110001001: DATA = 12'b011010001100;
            14'b00_111110001010: DATA = 12'b011010001111;
            14'b00_111110001011: DATA = 12'b011010010010;
            14'b00_111110001100: DATA = 12'b011010010101;
            14'b00_111110001101: DATA = 12'b011010011000;
            14'b00_111110001110: DATA = 12'b011010011011;
            14'b00_111110001111: DATA = 12'b011010011110;
            14'b00_111110010000: DATA = 12'b011010100010;
            14'b00_111110010001: DATA = 12'b011010100101;
            14'b00_111110010010: DATA = 12'b011010101000;
            14'b00_111110010011: DATA = 12'b011010101011;
            14'b00_111110010100: DATA = 12'b011010101110;
            14'b00_111110010101: DATA = 12'b011010110001;
            14'b00_111110010110: DATA = 12'b011010110100;
            14'b00_111110010111: DATA = 12'b011010110111;
            14'b00_111110011000: DATA = 12'b011010111010;
            14'b00_111110011001: DATA = 12'b011010111101;
            14'b00_111110011010: DATA = 12'b011011000001;
            14'b00_111110011011: DATA = 12'b011011000100;
            14'b00_111110011100: DATA = 12'b011011000111;
            14'b00_111110011101: DATA = 12'b011011001010;
            14'b00_111110011110: DATA = 12'b011011001101;
            14'b00_111110011111: DATA = 12'b011011010000;
            14'b00_111110100000: DATA = 12'b011011010011;
            14'b00_111110100001: DATA = 12'b011011010110;
            14'b00_111110100010: DATA = 12'b011011011001;
            14'b00_111110100011: DATA = 12'b011011011100;
            14'b00_111110100100: DATA = 12'b011011100000;
            14'b00_111110100101: DATA = 12'b011011100011;
            14'b00_111110100110: DATA = 12'b011011100110;
            14'b00_111110100111: DATA = 12'b011011101001;
            14'b00_111110101000: DATA = 12'b011011101100;
            14'b00_111110101001: DATA = 12'b011011101111;
            14'b00_111110101010: DATA = 12'b011011110010;
            14'b00_111110101011: DATA = 12'b011011110101;
            14'b00_111110101100: DATA = 12'b011011111000;
            14'b00_111110101101: DATA = 12'b011011111100;
            14'b00_111110101110: DATA = 12'b011011111111;
            14'b00_111110101111: DATA = 12'b011100000010;
            14'b00_111110110000: DATA = 12'b011100000101;
            14'b00_111110110001: DATA = 12'b011100001000;
            14'b00_111110110010: DATA = 12'b011100001011;
            14'b00_111110110011: DATA = 12'b011100001110;
            14'b00_111110110100: DATA = 12'b011100010001;
            14'b00_111110110101: DATA = 12'b011100010101;
            14'b00_111110110110: DATA = 12'b011100011000;
            14'b00_111110110111: DATA = 12'b011100011011;
            14'b00_111110111000: DATA = 12'b011100011110;
            14'b00_111110111001: DATA = 12'b011100100001;
            14'b00_111110111010: DATA = 12'b011100100100;
            14'b00_111110111011: DATA = 12'b011100100111;
            14'b00_111110111100: DATA = 12'b011100101010;
            14'b00_111110111101: DATA = 12'b011100101101;
            14'b00_111110111110: DATA = 12'b011100110001;
            14'b00_111110111111: DATA = 12'b011100110100;
            14'b00_111111000000: DATA = 12'b011100110111;
            14'b00_111111000001: DATA = 12'b011100111010;
            14'b00_111111000010: DATA = 12'b011100111101;
            14'b00_111111000011: DATA = 12'b011101000000;
            14'b00_111111000100: DATA = 12'b011101000011;
            14'b00_111111000101: DATA = 12'b011101000110;
            14'b00_111111000110: DATA = 12'b011101001010;
            14'b00_111111000111: DATA = 12'b011101001101;
            14'b00_111111001000: DATA = 12'b011101010000;
            14'b00_111111001001: DATA = 12'b011101010011;
            14'b00_111111001010: DATA = 12'b011101010110;
            14'b00_111111001011: DATA = 12'b011101011001;
            14'b00_111111001100: DATA = 12'b011101011100;
            14'b00_111111001101: DATA = 12'b011101100000;
            14'b00_111111001110: DATA = 12'b011101100011;
            14'b00_111111001111: DATA = 12'b011101100110;
            14'b00_111111010000: DATA = 12'b011101101001;
            14'b00_111111010001: DATA = 12'b011101101100;
            14'b00_111111010010: DATA = 12'b011101101111;
            14'b00_111111010011: DATA = 12'b011101110010;
            14'b00_111111010100: DATA = 12'b011101110101;
            14'b00_111111010101: DATA = 12'b011101111001;
            14'b00_111111010110: DATA = 12'b011101111100;
            14'b00_111111010111: DATA = 12'b011101111111;
            14'b00_111111011000: DATA = 12'b011110000010;
            14'b00_111111011001: DATA = 12'b011110000101;
            14'b00_111111011010: DATA = 12'b011110001000;
            14'b00_111111011011: DATA = 12'b011110001011;
            14'b00_111111011100: DATA = 12'b011110001111;
            14'b00_111111011101: DATA = 12'b011110010010;
            14'b00_111111011110: DATA = 12'b011110010101;
            14'b00_111111011111: DATA = 12'b011110011000;
            14'b00_111111100000: DATA = 12'b011110011011;
            14'b00_111111100001: DATA = 12'b011110011110;
            14'b00_111111100010: DATA = 12'b011110100001;
            14'b00_111111100011: DATA = 12'b011110100100;
            14'b00_111111100100: DATA = 12'b011110101000;
            14'b00_111111100101: DATA = 12'b011110101011;
            14'b00_111111100110: DATA = 12'b011110101110;
            14'b00_111111100111: DATA = 12'b011110110001;
            14'b00_111111101000: DATA = 12'b011110110100;
            14'b00_111111101001: DATA = 12'b011110110111;
            14'b00_111111101010: DATA = 12'b011110111010;
            14'b00_111111101011: DATA = 12'b011110111110;
            14'b00_111111101100: DATA = 12'b011111000001;
            14'b00_111111101101: DATA = 12'b011111000100;
            14'b00_111111101110: DATA = 12'b011111000111;
            14'b00_111111101111: DATA = 12'b011111001010;
            14'b00_111111110000: DATA = 12'b011111001101;
            14'b00_111111110001: DATA = 12'b011111010000;
            14'b00_111111110010: DATA = 12'b011111010100;
            14'b00_111111110011: DATA = 12'b011111010111;
            14'b00_111111110100: DATA = 12'b011111011010;
            14'b00_111111110101: DATA = 12'b011111011101;
            14'b00_111111110110: DATA = 12'b011111100000;
            14'b00_111111110111: DATA = 12'b011111100011;
            14'b00_111111111000: DATA = 12'b011111100110;
            14'b00_111111111001: DATA = 12'b011111101010;
            14'b00_111111111010: DATA = 12'b011111101101;
            14'b00_111111111011: DATA = 12'b011111110000;
            14'b00_111111111100: DATA = 12'b011111110011;
            14'b00_111111111101: DATA = 12'b011111110110;
            14'b00_111111111110: DATA = 12'b011111111001;
            14'b00_111111111111: DATA = 12'b011111111100;
            14'b01_000000000000: DATA = 12'b100000000000;
            14'b01_000000000001: DATA = 12'b100000000011;
            14'b01_000000000010: DATA = 12'b100000000110;
            14'b01_000000000011: DATA = 12'b100000001001;
            14'b01_000000000100: DATA = 12'b100000001100;
            14'b01_000000000101: DATA = 12'b100000001111;
            14'b01_000000000110: DATA = 12'b100000010010;
            14'b01_000000000111: DATA = 12'b100000010101;
            14'b01_000000001000: DATA = 12'b100000011001;
            14'b01_000000001001: DATA = 12'b100000011100;
            14'b01_000000001010: DATA = 12'b100000011111;
            14'b01_000000001011: DATA = 12'b100000100010;
            14'b01_000000001100: DATA = 12'b100000100101;
            14'b01_000000001101: DATA = 12'b100000101000;
            14'b01_000000001110: DATA = 12'b100000101011;
            14'b01_000000001111: DATA = 12'b100000101111;
            14'b01_000000010000: DATA = 12'b100000110010;
            14'b01_000000010001: DATA = 12'b100000110101;
            14'b01_000000010010: DATA = 12'b100000111000;
            14'b01_000000010011: DATA = 12'b100000111011;
            14'b01_000000010100: DATA = 12'b100000111110;
            14'b01_000000010101: DATA = 12'b100001000001;
            14'b01_000000010110: DATA = 12'b100001000101;
            14'b01_000000010111: DATA = 12'b100001001000;
            14'b01_000000011000: DATA = 12'b100001001011;
            14'b01_000000011001: DATA = 12'b100001001110;
            14'b01_000000011010: DATA = 12'b100001010001;
            14'b01_000000011011: DATA = 12'b100001010100;
            14'b01_000000011100: DATA = 12'b100001010111;
            14'b01_000000011101: DATA = 12'b100001011011;
            14'b01_000000011110: DATA = 12'b100001011110;
            14'b01_000000011111: DATA = 12'b100001100001;
            14'b01_000000100000: DATA = 12'b100001100100;
            14'b01_000000100001: DATA = 12'b100001100111;
            14'b01_000000100010: DATA = 12'b100001101010;
            14'b01_000000100011: DATA = 12'b100001101101;
            14'b01_000000100100: DATA = 12'b100001110000;
            14'b01_000000100101: DATA = 12'b100001110100;
            14'b01_000000100110: DATA = 12'b100001110111;
            14'b01_000000100111: DATA = 12'b100001111010;
            14'b01_000000101000: DATA = 12'b100001111101;
            14'b01_000000101001: DATA = 12'b100010000000;
            14'b01_000000101010: DATA = 12'b100010000011;
            14'b01_000000101011: DATA = 12'b100010000110;
            14'b01_000000101100: DATA = 12'b100010001010;
            14'b01_000000101101: DATA = 12'b100010001101;
            14'b01_000000101110: DATA = 12'b100010010000;
            14'b01_000000101111: DATA = 12'b100010010011;
            14'b01_000000110000: DATA = 12'b100010010110;
            14'b01_000000110001: DATA = 12'b100010011001;
            14'b01_000000110010: DATA = 12'b100010011100;
            14'b01_000000110011: DATA = 12'b100010011111;
            14'b01_000000110100: DATA = 12'b100010100011;
            14'b01_000000110101: DATA = 12'b100010100110;
            14'b01_000000110110: DATA = 12'b100010101001;
            14'b01_000000110111: DATA = 12'b100010101100;
            14'b01_000000111000: DATA = 12'b100010101111;
            14'b01_000000111001: DATA = 12'b100010110010;
            14'b01_000000111010: DATA = 12'b100010110101;
            14'b01_000000111011: DATA = 12'b100010111001;
            14'b01_000000111100: DATA = 12'b100010111100;
            14'b01_000000111101: DATA = 12'b100010111111;
            14'b01_000000111110: DATA = 12'b100011000010;
            14'b01_000000111111: DATA = 12'b100011000101;
            14'b01_000001000000: DATA = 12'b100011001000;
            14'b01_000001000001: DATA = 12'b100011001011;
            14'b01_000001000010: DATA = 12'b100011001110;
            14'b01_000001000011: DATA = 12'b100011010010;
            14'b01_000001000100: DATA = 12'b100011010101;
            14'b01_000001000101: DATA = 12'b100011011000;
            14'b01_000001000110: DATA = 12'b100011011011;
            14'b01_000001000111: DATA = 12'b100011011110;
            14'b01_000001001000: DATA = 12'b100011100001;
            14'b01_000001001001: DATA = 12'b100011100100;
            14'b01_000001001010: DATA = 12'b100011100111;
            14'b01_000001001011: DATA = 12'b100011101010;
            14'b01_000001001100: DATA = 12'b100011101110;
            14'b01_000001001101: DATA = 12'b100011110001;
            14'b01_000001001110: DATA = 12'b100011110100;
            14'b01_000001001111: DATA = 12'b100011110111;
            14'b01_000001010000: DATA = 12'b100011111010;
            14'b01_000001010001: DATA = 12'b100011111101;
            14'b01_000001010010: DATA = 12'b100100000000;
            14'b01_000001010011: DATA = 12'b100100000011;
            14'b01_000001010100: DATA = 12'b100100000111;
            14'b01_000001010101: DATA = 12'b100100001010;
            14'b01_000001010110: DATA = 12'b100100001101;
            14'b01_000001010111: DATA = 12'b100100010000;
            14'b01_000001011000: DATA = 12'b100100010011;
            14'b01_000001011001: DATA = 12'b100100010110;
            14'b01_000001011010: DATA = 12'b100100011001;
            14'b01_000001011011: DATA = 12'b100100011100;
            14'b01_000001011100: DATA = 12'b100100011111;
            14'b01_000001011101: DATA = 12'b100100100011;
            14'b01_000001011110: DATA = 12'b100100100110;
            14'b01_000001011111: DATA = 12'b100100101001;
            14'b01_000001100000: DATA = 12'b100100101100;
            14'b01_000001100001: DATA = 12'b100100101111;
            14'b01_000001100010: DATA = 12'b100100110010;
            14'b01_000001100011: DATA = 12'b100100110101;
            14'b01_000001100100: DATA = 12'b100100111000;
            14'b01_000001100101: DATA = 12'b100100111011;
            14'b01_000001100110: DATA = 12'b100100111110;
            14'b01_000001100111: DATA = 12'b100101000010;
            14'b01_000001101000: DATA = 12'b100101000101;
            14'b01_000001101001: DATA = 12'b100101001000;
            14'b01_000001101010: DATA = 12'b100101001011;
            14'b01_000001101011: DATA = 12'b100101001110;
            14'b01_000001101100: DATA = 12'b100101010001;
            14'b01_000001101101: DATA = 12'b100101010100;
            14'b01_000001101110: DATA = 12'b100101010111;
            14'b01_000001101111: DATA = 12'b100101011010;
            14'b01_000001110000: DATA = 12'b100101011101;
            14'b01_000001110001: DATA = 12'b100101100001;
            14'b01_000001110010: DATA = 12'b100101100100;
            14'b01_000001110011: DATA = 12'b100101100111;
            14'b01_000001110100: DATA = 12'b100101101010;
            14'b01_000001110101: DATA = 12'b100101101101;
            14'b01_000001110110: DATA = 12'b100101110000;
            14'b01_000001110111: DATA = 12'b100101110011;
            14'b01_000001111000: DATA = 12'b100101110110;
            14'b01_000001111001: DATA = 12'b100101111001;
            14'b01_000001111010: DATA = 12'b100101111100;
            14'b01_000001111011: DATA = 12'b100101111111;
            14'b01_000001111100: DATA = 12'b100110000011;
            14'b01_000001111101: DATA = 12'b100110000110;
            14'b01_000001111110: DATA = 12'b100110001001;
            14'b01_000001111111: DATA = 12'b100110001100;
            14'b01_000010000000: DATA = 12'b100110001111;
            14'b01_000010000001: DATA = 12'b100110010010;
            14'b01_000010000010: DATA = 12'b100110010101;
            14'b01_000010000011: DATA = 12'b100110011000;
            14'b01_000010000100: DATA = 12'b100110011011;
            14'b01_000010000101: DATA = 12'b100110011110;
            14'b01_000010000110: DATA = 12'b100110100001;
            14'b01_000010000111: DATA = 12'b100110100100;
            14'b01_000010001000: DATA = 12'b100110100111;
            14'b01_000010001001: DATA = 12'b100110101011;
            14'b01_000010001010: DATA = 12'b100110101110;
            14'b01_000010001011: DATA = 12'b100110110001;
            14'b01_000010001100: DATA = 12'b100110110100;
            14'b01_000010001101: DATA = 12'b100110110111;
            14'b01_000010001110: DATA = 12'b100110111010;
            14'b01_000010001111: DATA = 12'b100110111101;
            14'b01_000010010000: DATA = 12'b100111000000;
            14'b01_000010010001: DATA = 12'b100111000011;
            14'b01_000010010010: DATA = 12'b100111000110;
            14'b01_000010010011: DATA = 12'b100111001001;
            14'b01_000010010100: DATA = 12'b100111001100;
            14'b01_000010010101: DATA = 12'b100111001111;
            14'b01_000010010110: DATA = 12'b100111010010;
            14'b01_000010010111: DATA = 12'b100111010101;
            14'b01_000010011000: DATA = 12'b100111011000;
            14'b01_000010011001: DATA = 12'b100111011100;
            14'b01_000010011010: DATA = 12'b100111011111;
            14'b01_000010011011: DATA = 12'b100111100010;
            14'b01_000010011100: DATA = 12'b100111100101;
            14'b01_000010011101: DATA = 12'b100111101000;
            14'b01_000010011110: DATA = 12'b100111101011;
            14'b01_000010011111: DATA = 12'b100111101110;
            14'b01_000010100000: DATA = 12'b100111110001;
            14'b01_000010100001: DATA = 12'b100111110100;
            14'b01_000010100010: DATA = 12'b100111110111;
            14'b01_000010100011: DATA = 12'b100111111010;
            14'b01_000010100100: DATA = 12'b100111111101;
            14'b01_000010100101: DATA = 12'b101000000000;
            14'b01_000010100110: DATA = 12'b101000000011;
            14'b01_000010100111: DATA = 12'b101000000110;
            14'b01_000010101000: DATA = 12'b101000001001;
            14'b01_000010101001: DATA = 12'b101000001100;
            14'b01_000010101010: DATA = 12'b101000001111;
            14'b01_000010101011: DATA = 12'b101000010010;
            14'b01_000010101100: DATA = 12'b101000010101;
            14'b01_000010101101: DATA = 12'b101000011000;
            14'b01_000010101110: DATA = 12'b101000011011;
            14'b01_000010101111: DATA = 12'b101000011110;
            14'b01_000010110000: DATA = 12'b101000100001;
            14'b01_000010110001: DATA = 12'b101000100100;
            14'b01_000010110010: DATA = 12'b101000101000;
            14'b01_000010110011: DATA = 12'b101000101011;
            14'b01_000010110100: DATA = 12'b101000101110;
            14'b01_000010110101: DATA = 12'b101000110001;
            14'b01_000010110110: DATA = 12'b101000110100;
            14'b01_000010110111: DATA = 12'b101000110111;
            14'b01_000010111000: DATA = 12'b101000111010;
            14'b01_000010111001: DATA = 12'b101000111101;
            14'b01_000010111010: DATA = 12'b101001000000;
            14'b01_000010111011: DATA = 12'b101001000011;
            14'b01_000010111100: DATA = 12'b101001000110;
            14'b01_000010111101: DATA = 12'b101001001001;
            14'b01_000010111110: DATA = 12'b101001001100;
            14'b01_000010111111: DATA = 12'b101001001111;
            14'b01_000011000000: DATA = 12'b101001010010;
            14'b01_000011000001: DATA = 12'b101001010101;
            14'b01_000011000010: DATA = 12'b101001011000;
            14'b01_000011000011: DATA = 12'b101001011011;
            14'b01_000011000100: DATA = 12'b101001011110;
            14'b01_000011000101: DATA = 12'b101001100001;
            14'b01_000011000110: DATA = 12'b101001100100;
            14'b01_000011000111: DATA = 12'b101001100111;
            14'b01_000011001000: DATA = 12'b101001101010;
            14'b01_000011001001: DATA = 12'b101001101101;
            14'b01_000011001010: DATA = 12'b101001110000;
            14'b01_000011001011: DATA = 12'b101001110011;
            14'b01_000011001100: DATA = 12'b101001110110;
            14'b01_000011001101: DATA = 12'b101001111001;
            14'b01_000011001110: DATA = 12'b101001111100;
            14'b01_000011001111: DATA = 12'b101001111111;
            14'b01_000011010000: DATA = 12'b101010000010;
            14'b01_000011010001: DATA = 12'b101010000101;
            14'b01_000011010010: DATA = 12'b101010001000;
            14'b01_000011010011: DATA = 12'b101010001011;
            14'b01_000011010100: DATA = 12'b101010001110;
            14'b01_000011010101: DATA = 12'b101010010000;
            14'b01_000011010110: DATA = 12'b101010010011;
            14'b01_000011010111: DATA = 12'b101010010110;
            14'b01_000011011000: DATA = 12'b101010011001;
            14'b01_000011011001: DATA = 12'b101010011100;
            14'b01_000011011010: DATA = 12'b101010011111;
            14'b01_000011011011: DATA = 12'b101010100010;
            14'b01_000011011100: DATA = 12'b101010100101;
            14'b01_000011011101: DATA = 12'b101010101000;
            14'b01_000011011110: DATA = 12'b101010101011;
            14'b01_000011011111: DATA = 12'b101010101110;
            14'b01_000011100000: DATA = 12'b101010110001;
            14'b01_000011100001: DATA = 12'b101010110100;
            14'b01_000011100010: DATA = 12'b101010110111;
            14'b01_000011100011: DATA = 12'b101010111010;
            14'b01_000011100100: DATA = 12'b101010111101;
            14'b01_000011100101: DATA = 12'b101011000000;
            14'b01_000011100110: DATA = 12'b101011000011;
            14'b01_000011100111: DATA = 12'b101011000110;
            14'b01_000011101000: DATA = 12'b101011001001;
            14'b01_000011101001: DATA = 12'b101011001100;
            14'b01_000011101010: DATA = 12'b101011001111;
            14'b01_000011101011: DATA = 12'b101011010010;
            14'b01_000011101100: DATA = 12'b101011010100;
            14'b01_000011101101: DATA = 12'b101011010111;
            14'b01_000011101110: DATA = 12'b101011011010;
            14'b01_000011101111: DATA = 12'b101011011101;
            14'b01_000011110000: DATA = 12'b101011100000;
            14'b01_000011110001: DATA = 12'b101011100011;
            14'b01_000011110010: DATA = 12'b101011100110;
            14'b01_000011110011: DATA = 12'b101011101001;
            14'b01_000011110100: DATA = 12'b101011101100;
            14'b01_000011110101: DATA = 12'b101011101111;
            14'b01_000011110110: DATA = 12'b101011110010;
            14'b01_000011110111: DATA = 12'b101011110101;
            14'b01_000011111000: DATA = 12'b101011111000;
            14'b01_000011111001: DATA = 12'b101011111011;
            14'b01_000011111010: DATA = 12'b101011111101;
            14'b01_000011111011: DATA = 12'b101100000000;
            14'b01_000011111100: DATA = 12'b101100000011;
            14'b01_000011111101: DATA = 12'b101100000110;
            14'b01_000011111110: DATA = 12'b101100001001;
            14'b01_000011111111: DATA = 12'b101100001100;
            14'b01_000100000000: DATA = 12'b101100001111;
            14'b01_000100000001: DATA = 12'b101100010010;
            14'b01_000100000010: DATA = 12'b101100010101;
            14'b01_000100000011: DATA = 12'b101100011000;
            14'b01_000100000100: DATA = 12'b101100011010;
            14'b01_000100000101: DATA = 12'b101100011101;
            14'b01_000100000110: DATA = 12'b101100100000;
            14'b01_000100000111: DATA = 12'b101100100011;
            14'b01_000100001000: DATA = 12'b101100100110;
            14'b01_000100001001: DATA = 12'b101100101001;
            14'b01_000100001010: DATA = 12'b101100101100;
            14'b01_000100001011: DATA = 12'b101100101111;
            14'b01_000100001100: DATA = 12'b101100110010;
            14'b01_000100001101: DATA = 12'b101100110100;
            14'b01_000100001110: DATA = 12'b101100110111;
            14'b01_000100001111: DATA = 12'b101100111010;
            14'b01_000100010000: DATA = 12'b101100111101;
            14'b01_000100010001: DATA = 12'b101101000000;
            14'b01_000100010010: DATA = 12'b101101000011;
            14'b01_000100010011: DATA = 12'b101101000110;
            14'b01_000100010100: DATA = 12'b101101001000;
            14'b01_000100010101: DATA = 12'b101101001011;
            14'b01_000100010110: DATA = 12'b101101001110;
            14'b01_000100010111: DATA = 12'b101101010001;
            14'b01_000100011000: DATA = 12'b101101010100;
            14'b01_000100011001: DATA = 12'b101101010111;
            14'b01_000100011010: DATA = 12'b101101011010;
            14'b01_000100011011: DATA = 12'b101101011100;
            14'b01_000100011100: DATA = 12'b101101011111;
            14'b01_000100011101: DATA = 12'b101101100010;
            14'b01_000100011110: DATA = 12'b101101100101;
            14'b01_000100011111: DATA = 12'b101101101000;
            14'b01_000100100000: DATA = 12'b101101101011;
            14'b01_000100100001: DATA = 12'b101101101110;
            14'b01_000100100010: DATA = 12'b101101110000;
            14'b01_000100100011: DATA = 12'b101101110011;
            14'b01_000100100100: DATA = 12'b101101110110;
            14'b01_000100100101: DATA = 12'b101101111001;
            14'b01_000100100110: DATA = 12'b101101111100;
            14'b01_000100100111: DATA = 12'b101101111111;
            14'b01_000100101000: DATA = 12'b101110000001;
            14'b01_000100101001: DATA = 12'b101110000100;
            14'b01_000100101010: DATA = 12'b101110000111;
            14'b01_000100101011: DATA = 12'b101110001010;
            14'b01_000100101100: DATA = 12'b101110001101;
            14'b01_000100101101: DATA = 12'b101110001111;
            14'b01_000100101110: DATA = 12'b101110010010;
            14'b01_000100101111: DATA = 12'b101110010101;
            14'b01_000100110000: DATA = 12'b101110011000;
            14'b01_000100110001: DATA = 12'b101110011011;
            14'b01_000100110010: DATA = 12'b101110011101;
            14'b01_000100110011: DATA = 12'b101110100000;
            14'b01_000100110100: DATA = 12'b101110100011;
            14'b01_000100110101: DATA = 12'b101110100110;
            14'b01_000100110110: DATA = 12'b101110101001;
            14'b01_000100110111: DATA = 12'b101110101011;
            14'b01_000100111000: DATA = 12'b101110101110;
            14'b01_000100111001: DATA = 12'b101110110001;
            14'b01_000100111010: DATA = 12'b101110110100;
            14'b01_000100111011: DATA = 12'b101110110111;
            14'b01_000100111100: DATA = 12'b101110111001;
            14'b01_000100111101: DATA = 12'b101110111100;
            14'b01_000100111110: DATA = 12'b101110111111;
            14'b01_000100111111: DATA = 12'b101111000010;
            14'b01_000101000000: DATA = 12'b101111000100;
            14'b01_000101000001: DATA = 12'b101111000111;
            14'b01_000101000010: DATA = 12'b101111001010;
            14'b01_000101000011: DATA = 12'b101111001101;
            14'b01_000101000100: DATA = 12'b101111010000;
            14'b01_000101000101: DATA = 12'b101111010010;
            14'b01_000101000110: DATA = 12'b101111010101;
            14'b01_000101000111: DATA = 12'b101111011000;
            14'b01_000101001000: DATA = 12'b101111011011;
            14'b01_000101001001: DATA = 12'b101111011101;
            14'b01_000101001010: DATA = 12'b101111100000;
            14'b01_000101001011: DATA = 12'b101111100011;
            14'b01_000101001100: DATA = 12'b101111100110;
            14'b01_000101001101: DATA = 12'b101111101000;
            14'b01_000101001110: DATA = 12'b101111101011;
            14'b01_000101001111: DATA = 12'b101111101110;
            14'b01_000101010000: DATA = 12'b101111110000;
            14'b01_000101010001: DATA = 12'b101111110011;
            14'b01_000101010010: DATA = 12'b101111110110;
            14'b01_000101010011: DATA = 12'b101111111001;
            14'b01_000101010100: DATA = 12'b101111111011;
            14'b01_000101010101: DATA = 12'b101111111110;
            14'b01_000101010110: DATA = 12'b110000000001;
            14'b01_000101010111: DATA = 12'b110000000100;
            14'b01_000101011000: DATA = 12'b110000000110;
            14'b01_000101011001: DATA = 12'b110000001001;
            14'b01_000101011010: DATA = 12'b110000001100;
            14'b01_000101011011: DATA = 12'b110000001110;
            14'b01_000101011100: DATA = 12'b110000010001;
            14'b01_000101011101: DATA = 12'b110000010100;
            14'b01_000101011110: DATA = 12'b110000010110;
            14'b01_000101011111: DATA = 12'b110000011001;
            14'b01_000101100000: DATA = 12'b110000011100;
            14'b01_000101100001: DATA = 12'b110000011111;
            14'b01_000101100010: DATA = 12'b110000100001;
            14'b01_000101100011: DATA = 12'b110000100100;
            14'b01_000101100100: DATA = 12'b110000100111;
            14'b01_000101100101: DATA = 12'b110000101001;
            14'b01_000101100110: DATA = 12'b110000101100;
            14'b01_000101100111: DATA = 12'b110000101111;
            14'b01_000101101000: DATA = 12'b110000110001;
            14'b01_000101101001: DATA = 12'b110000110100;
            14'b01_000101101010: DATA = 12'b110000110111;
            14'b01_000101101011: DATA = 12'b110000111001;
            14'b01_000101101100: DATA = 12'b110000111100;
            14'b01_000101101101: DATA = 12'b110000111111;
            14'b01_000101101110: DATA = 12'b110001000001;
            14'b01_000101101111: DATA = 12'b110001000100;
            14'b01_000101110000: DATA = 12'b110001000111;
            14'b01_000101110001: DATA = 12'b110001001001;
            14'b01_000101110010: DATA = 12'b110001001100;
            14'b01_000101110011: DATA = 12'b110001001111;
            14'b01_000101110100: DATA = 12'b110001010001;
            14'b01_000101110101: DATA = 12'b110001010100;
            14'b01_000101110110: DATA = 12'b110001010111;
            14'b01_000101110111: DATA = 12'b110001011001;
            14'b01_000101111000: DATA = 12'b110001011100;
            14'b01_000101111001: DATA = 12'b110001011110;
            14'b01_000101111010: DATA = 12'b110001100001;
            14'b01_000101111011: DATA = 12'b110001100100;
            14'b01_000101111100: DATA = 12'b110001100110;
            14'b01_000101111101: DATA = 12'b110001101001;
            14'b01_000101111110: DATA = 12'b110001101100;
            14'b01_000101111111: DATA = 12'b110001101110;
            14'b01_000110000000: DATA = 12'b110001110001;
            14'b01_000110000001: DATA = 12'b110001110011;
            14'b01_000110000010: DATA = 12'b110001110110;
            14'b01_000110000011: DATA = 12'b110001111001;
            14'b01_000110000100: DATA = 12'b110001111011;
            14'b01_000110000101: DATA = 12'b110001111110;
            14'b01_000110000110: DATA = 12'b110010000000;
            14'b01_000110000111: DATA = 12'b110010000011;
            14'b01_000110001000: DATA = 12'b110010000110;
            14'b01_000110001001: DATA = 12'b110010001000;
            14'b01_000110001010: DATA = 12'b110010001011;
            14'b01_000110001011: DATA = 12'b110010001101;
            14'b01_000110001100: DATA = 12'b110010010000;
            14'b01_000110001101: DATA = 12'b110010010010;
            14'b01_000110001110: DATA = 12'b110010010101;
            14'b01_000110001111: DATA = 12'b110010011000;
            14'b01_000110010000: DATA = 12'b110010011010;
            14'b01_000110010001: DATA = 12'b110010011101;
            14'b01_000110010010: DATA = 12'b110010011111;
            14'b01_000110010011: DATA = 12'b110010100010;
            14'b01_000110010100: DATA = 12'b110010100100;
            14'b01_000110010101: DATA = 12'b110010100111;
            14'b01_000110010110: DATA = 12'b110010101010;
            14'b01_000110010111: DATA = 12'b110010101100;
            14'b01_000110011000: DATA = 12'b110010101111;
            14'b01_000110011001: DATA = 12'b110010110001;
            14'b01_000110011010: DATA = 12'b110010110100;
            14'b01_000110011011: DATA = 12'b110010110110;
            14'b01_000110011100: DATA = 12'b110010111001;
            14'b01_000110011101: DATA = 12'b110010111011;
            14'b01_000110011110: DATA = 12'b110010111110;
            14'b01_000110011111: DATA = 12'b110011000000;
            14'b01_000110100000: DATA = 12'b110011000011;
            14'b01_000110100001: DATA = 12'b110011000101;
            14'b01_000110100010: DATA = 12'b110011001000;
            14'b01_000110100011: DATA = 12'b110011001010;
            14'b01_000110100100: DATA = 12'b110011001101;
            14'b01_000110100101: DATA = 12'b110011001111;
            14'b01_000110100110: DATA = 12'b110011010010;
            14'b01_000110100111: DATA = 12'b110011010100;
            14'b01_000110101000: DATA = 12'b110011010111;
            14'b01_000110101001: DATA = 12'b110011011001;
            14'b01_000110101010: DATA = 12'b110011011100;
            14'b01_000110101011: DATA = 12'b110011011110;
            14'b01_000110101100: DATA = 12'b110011100001;
            14'b01_000110101101: DATA = 12'b110011100011;
            14'b01_000110101110: DATA = 12'b110011100110;
            14'b01_000110101111: DATA = 12'b110011101000;
            14'b01_000110110000: DATA = 12'b110011101011;
            14'b01_000110110001: DATA = 12'b110011101101;
            14'b01_000110110010: DATA = 12'b110011110000;
            14'b01_000110110011: DATA = 12'b110011110010;
            14'b01_000110110100: DATA = 12'b110011110101;
            14'b01_000110110101: DATA = 12'b110011110111;
            14'b01_000110110110: DATA = 12'b110011111010;
            14'b01_000110110111: DATA = 12'b110011111100;
            14'b01_000110111000: DATA = 12'b110011111111;
            14'b01_000110111001: DATA = 12'b110100000001;
            14'b01_000110111010: DATA = 12'b110100000011;
            14'b01_000110111011: DATA = 12'b110100000110;
            14'b01_000110111100: DATA = 12'b110100001000;
            14'b01_000110111101: DATA = 12'b110100001011;
            14'b01_000110111110: DATA = 12'b110100001101;
            14'b01_000110111111: DATA = 12'b110100010000;
            14'b01_000111000000: DATA = 12'b110100010010;
            14'b01_000111000001: DATA = 12'b110100010101;
            14'b01_000111000010: DATA = 12'b110100010111;
            14'b01_000111000011: DATA = 12'b110100011001;
            14'b01_000111000100: DATA = 12'b110100011100;
            14'b01_000111000101: DATA = 12'b110100011110;
            14'b01_000111000110: DATA = 12'b110100100001;
            14'b01_000111000111: DATA = 12'b110100100011;
            14'b01_000111001000: DATA = 12'b110100100101;
            14'b01_000111001001: DATA = 12'b110100101000;
            14'b01_000111001010: DATA = 12'b110100101010;
            14'b01_000111001011: DATA = 12'b110100101101;
            14'b01_000111001100: DATA = 12'b110100101111;
            14'b01_000111001101: DATA = 12'b110100110001;
            14'b01_000111001110: DATA = 12'b110100110100;
            14'b01_000111001111: DATA = 12'b110100110110;
            14'b01_000111010000: DATA = 12'b110100111001;
            14'b01_000111010001: DATA = 12'b110100111011;
            14'b01_000111010010: DATA = 12'b110100111101;
            14'b01_000111010011: DATA = 12'b110101000000;
            14'b01_000111010100: DATA = 12'b110101000010;
            14'b01_000111010101: DATA = 12'b110101000100;
            14'b01_000111010110: DATA = 12'b110101000111;
            14'b01_000111010111: DATA = 12'b110101001001;
            14'b01_000111011000: DATA = 12'b110101001011;
            14'b01_000111011001: DATA = 12'b110101001110;
            14'b01_000111011010: DATA = 12'b110101010000;
            14'b01_000111011011: DATA = 12'b110101010011;
            14'b01_000111011100: DATA = 12'b110101010101;
            14'b01_000111011101: DATA = 12'b110101010111;
            14'b01_000111011110: DATA = 12'b110101011010;
            14'b01_000111011111: DATA = 12'b110101011100;
            14'b01_000111100000: DATA = 12'b110101011110;
            14'b01_000111100001: DATA = 12'b110101100001;
            14'b01_000111100010: DATA = 12'b110101100011;
            14'b01_000111100011: DATA = 12'b110101100101;
            14'b01_000111100100: DATA = 12'b110101100111;
            14'b01_000111100101: DATA = 12'b110101101010;
            14'b01_000111100110: DATA = 12'b110101101100;
            14'b01_000111100111: DATA = 12'b110101101110;
            14'b01_000111101000: DATA = 12'b110101110001;
            14'b01_000111101001: DATA = 12'b110101110011;
            14'b01_000111101010: DATA = 12'b110101110101;
            14'b01_000111101011: DATA = 12'b110101111000;
            14'b01_000111101100: DATA = 12'b110101111010;
            14'b01_000111101101: DATA = 12'b110101111100;
            14'b01_000111101110: DATA = 12'b110101111110;
            14'b01_000111101111: DATA = 12'b110110000001;
            14'b01_000111110000: DATA = 12'b110110000011;
            14'b01_000111110001: DATA = 12'b110110000101;
            14'b01_000111110010: DATA = 12'b110110001000;
            14'b01_000111110011: DATA = 12'b110110001010;
            14'b01_000111110100: DATA = 12'b110110001100;
            14'b01_000111110101: DATA = 12'b110110001110;
            14'b01_000111110110: DATA = 12'b110110010001;
            14'b01_000111110111: DATA = 12'b110110010011;
            14'b01_000111111000: DATA = 12'b110110010101;
            14'b01_000111111001: DATA = 12'b110110010111;
            14'b01_000111111010: DATA = 12'b110110011010;
            14'b01_000111111011: DATA = 12'b110110011100;
            14'b01_000111111100: DATA = 12'b110110011110;
            14'b01_000111111101: DATA = 12'b110110100000;
            14'b01_000111111110: DATA = 12'b110110100011;
            14'b01_000111111111: DATA = 12'b110110100101;
            14'b01_001000000000: DATA = 12'b110110100111;
            14'b01_001000000001: DATA = 12'b110110101001;
            14'b01_001000000010: DATA = 12'b110110101011;
            14'b01_001000000011: DATA = 12'b110110101110;
            14'b01_001000000100: DATA = 12'b110110110000;
            14'b01_001000000101: DATA = 12'b110110110010;
            14'b01_001000000110: DATA = 12'b110110110100;
            14'b01_001000000111: DATA = 12'b110110110110;
            14'b01_001000001000: DATA = 12'b110110111001;
            14'b01_001000001001: DATA = 12'b110110111011;
            14'b01_001000001010: DATA = 12'b110110111101;
            14'b01_001000001011: DATA = 12'b110110111111;
            14'b01_001000001100: DATA = 12'b110111000001;
            14'b01_001000001101: DATA = 12'b110111000100;
            14'b01_001000001110: DATA = 12'b110111000110;
            14'b01_001000001111: DATA = 12'b110111001000;
            14'b01_001000010000: DATA = 12'b110111001010;
            14'b01_001000010001: DATA = 12'b110111001100;
            14'b01_001000010010: DATA = 12'b110111001110;
            14'b01_001000010011: DATA = 12'b110111010001;
            14'b01_001000010100: DATA = 12'b110111010011;
            14'b01_001000010101: DATA = 12'b110111010101;
            14'b01_001000010110: DATA = 12'b110111010111;
            14'b01_001000010111: DATA = 12'b110111011001;
            14'b01_001000011000: DATA = 12'b110111011011;
            14'b01_001000011001: DATA = 12'b110111011101;
            14'b01_001000011010: DATA = 12'b110111100000;
            14'b01_001000011011: DATA = 12'b110111100010;
            14'b01_001000011100: DATA = 12'b110111100100;
            14'b01_001000011101: DATA = 12'b110111100110;
            14'b01_001000011110: DATA = 12'b110111101000;
            14'b01_001000011111: DATA = 12'b110111101010;
            14'b01_001000100000: DATA = 12'b110111101100;
            14'b01_001000100001: DATA = 12'b110111101110;
            14'b01_001000100010: DATA = 12'b110111110000;
            14'b01_001000100011: DATA = 12'b110111110011;
            14'b01_001000100100: DATA = 12'b110111110101;
            14'b01_001000100101: DATA = 12'b110111110111;
            14'b01_001000100110: DATA = 12'b110111111001;
            14'b01_001000100111: DATA = 12'b110111111011;
            14'b01_001000101000: DATA = 12'b110111111101;
            14'b01_001000101001: DATA = 12'b110111111111;
            14'b01_001000101010: DATA = 12'b111000000001;
            14'b01_001000101011: DATA = 12'b111000000011;
            14'b01_001000101100: DATA = 12'b111000000101;
            14'b01_001000101101: DATA = 12'b111000000111;
            14'b01_001000101110: DATA = 12'b111000001001;
            14'b01_001000101111: DATA = 12'b111000001011;
            14'b01_001000110000: DATA = 12'b111000001110;
            14'b01_001000110001: DATA = 12'b111000010000;
            14'b01_001000110010: DATA = 12'b111000010010;
            14'b01_001000110011: DATA = 12'b111000010100;
            14'b01_001000110100: DATA = 12'b111000010110;
            14'b01_001000110101: DATA = 12'b111000011000;
            14'b01_001000110110: DATA = 12'b111000011010;
            14'b01_001000110111: DATA = 12'b111000011100;
            14'b01_001000111000: DATA = 12'b111000011110;
            14'b01_001000111001: DATA = 12'b111000100000;
            14'b01_001000111010: DATA = 12'b111000100010;
            14'b01_001000111011: DATA = 12'b111000100100;
            14'b01_001000111100: DATA = 12'b111000100110;
            14'b01_001000111101: DATA = 12'b111000101000;
            14'b01_001000111110: DATA = 12'b111000101010;
            14'b01_001000111111: DATA = 12'b111000101100;
            14'b01_001001000000: DATA = 12'b111000101110;
            14'b01_001001000001: DATA = 12'b111000110000;
            14'b01_001001000010: DATA = 12'b111000110010;
            14'b01_001001000011: DATA = 12'b111000110100;
            14'b01_001001000100: DATA = 12'b111000110110;
            14'b01_001001000101: DATA = 12'b111000111000;
            14'b01_001001000110: DATA = 12'b111000111010;
            14'b01_001001000111: DATA = 12'b111000111100;
            14'b01_001001001000: DATA = 12'b111000111110;
            14'b01_001001001001: DATA = 12'b111001000000;
            14'b01_001001001010: DATA = 12'b111001000010;
            14'b01_001001001011: DATA = 12'b111001000100;
            14'b01_001001001100: DATA = 12'b111001000101;
            14'b01_001001001101: DATA = 12'b111001000111;
            14'b01_001001001110: DATA = 12'b111001001001;
            14'b01_001001001111: DATA = 12'b111001001011;
            14'b01_001001010000: DATA = 12'b111001001101;
            14'b01_001001010001: DATA = 12'b111001001111;
            14'b01_001001010010: DATA = 12'b111001010001;
            14'b01_001001010011: DATA = 12'b111001010011;
            14'b01_001001010100: DATA = 12'b111001010101;
            14'b01_001001010101: DATA = 12'b111001010111;
            14'b01_001001010110: DATA = 12'b111001011001;
            14'b01_001001010111: DATA = 12'b111001011011;
            14'b01_001001011000: DATA = 12'b111001011101;
            14'b01_001001011001: DATA = 12'b111001011110;
            14'b01_001001011010: DATA = 12'b111001100000;
            14'b01_001001011011: DATA = 12'b111001100010;
            14'b01_001001011100: DATA = 12'b111001100100;
            14'b01_001001011101: DATA = 12'b111001100110;
            14'b01_001001011110: DATA = 12'b111001101000;
            14'b01_001001011111: DATA = 12'b111001101010;
            14'b01_001001100000: DATA = 12'b111001101100;
            14'b01_001001100001: DATA = 12'b111001101110;
            14'b01_001001100010: DATA = 12'b111001101111;
            14'b01_001001100011: DATA = 12'b111001110001;
            14'b01_001001100100: DATA = 12'b111001110011;
            14'b01_001001100101: DATA = 12'b111001110101;
            14'b01_001001100110: DATA = 12'b111001110111;
            14'b01_001001100111: DATA = 12'b111001111001;
            14'b01_001001101000: DATA = 12'b111001111011;
            14'b01_001001101001: DATA = 12'b111001111100;
            14'b01_001001101010: DATA = 12'b111001111110;
            14'b01_001001101011: DATA = 12'b111010000000;
            14'b01_001001101100: DATA = 12'b111010000010;
            14'b01_001001101101: DATA = 12'b111010000100;
            14'b01_001001101110: DATA = 12'b111010000101;
            14'b01_001001101111: DATA = 12'b111010000111;
            14'b01_001001110000: DATA = 12'b111010001001;
            14'b01_001001110001: DATA = 12'b111010001011;
            14'b01_001001110010: DATA = 12'b111010001101;
            14'b01_001001110011: DATA = 12'b111010001111;
            14'b01_001001110100: DATA = 12'b111010010000;
            14'b01_001001110101: DATA = 12'b111010010010;
            14'b01_001001110110: DATA = 12'b111010010100;
            14'b01_001001110111: DATA = 12'b111010010110;
            14'b01_001001111000: DATA = 12'b111010010111;
            14'b01_001001111001: DATA = 12'b111010011001;
            14'b01_001001111010: DATA = 12'b111010011011;
            14'b01_001001111011: DATA = 12'b111010011101;
            14'b01_001001111100: DATA = 12'b111010011111;
            14'b01_001001111101: DATA = 12'b111010100000;
            14'b01_001001111110: DATA = 12'b111010100010;
            14'b01_001001111111: DATA = 12'b111010100100;
            14'b01_001010000000: DATA = 12'b111010100110;
            14'b01_001010000001: DATA = 12'b111010100111;
            14'b01_001010000010: DATA = 12'b111010101001;
            14'b01_001010000011: DATA = 12'b111010101011;
            14'b01_001010000100: DATA = 12'b111010101100;
            14'b01_001010000101: DATA = 12'b111010101110;
            14'b01_001010000110: DATA = 12'b111010110000;
            14'b01_001010000111: DATA = 12'b111010110010;
            14'b01_001010001000: DATA = 12'b111010110011;
            14'b01_001010001001: DATA = 12'b111010110101;
            14'b01_001010001010: DATA = 12'b111010110111;
            14'b01_001010001011: DATA = 12'b111010111000;
            14'b01_001010001100: DATA = 12'b111010111010;
            14'b01_001010001101: DATA = 12'b111010111100;
            14'b01_001010001110: DATA = 12'b111010111110;
            14'b01_001010001111: DATA = 12'b111010111111;
            14'b01_001010010000: DATA = 12'b111011000001;
            14'b01_001010010001: DATA = 12'b111011000011;
            14'b01_001010010010: DATA = 12'b111011000100;
            14'b01_001010010011: DATA = 12'b111011000110;
            14'b01_001010010100: DATA = 12'b111011001000;
            14'b01_001010010101: DATA = 12'b111011001001;
            14'b01_001010010110: DATA = 12'b111011001011;
            14'b01_001010010111: DATA = 12'b111011001101;
            14'b01_001010011000: DATA = 12'b111011001110;
            14'b01_001010011001: DATA = 12'b111011010000;
            14'b01_001010011010: DATA = 12'b111011010010;
            14'b01_001010011011: DATA = 12'b111011010011;
            14'b01_001010011100: DATA = 12'b111011010101;
            14'b01_001010011101: DATA = 12'b111011010110;
            14'b01_001010011110: DATA = 12'b111011011000;
            14'b01_001010011111: DATA = 12'b111011011010;
            14'b01_001010100000: DATA = 12'b111011011011;
            14'b01_001010100001: DATA = 12'b111011011101;
            14'b01_001010100010: DATA = 12'b111011011110;
            14'b01_001010100011: DATA = 12'b111011100000;
            14'b01_001010100100: DATA = 12'b111011100010;
            14'b01_001010100101: DATA = 12'b111011100011;
            14'b01_001010100110: DATA = 12'b111011100101;
            14'b01_001010100111: DATA = 12'b111011100110;
            14'b01_001010101000: DATA = 12'b111011101000;
            14'b01_001010101001: DATA = 12'b111011101010;
            14'b01_001010101010: DATA = 12'b111011101011;
            14'b01_001010101011: DATA = 12'b111011101101;
            14'b01_001010101100: DATA = 12'b111011101110;
            14'b01_001010101101: DATA = 12'b111011110000;
            14'b01_001010101110: DATA = 12'b111011110001;
            14'b01_001010101111: DATA = 12'b111011110011;
            14'b01_001010110000: DATA = 12'b111011110101;
            14'b01_001010110001: DATA = 12'b111011110110;
            14'b01_001010110010: DATA = 12'b111011111000;
            14'b01_001010110011: DATA = 12'b111011111001;
            14'b01_001010110100: DATA = 12'b111011111011;
            14'b01_001010110101: DATA = 12'b111011111100;
            14'b01_001010110110: DATA = 12'b111011111110;
            14'b01_001010110111: DATA = 12'b111011111111;
            14'b01_001010111000: DATA = 12'b111100000001;
            14'b01_001010111001: DATA = 12'b111100000010;
            14'b01_001010111010: DATA = 12'b111100000100;
            14'b01_001010111011: DATA = 12'b111100000101;
            14'b01_001010111100: DATA = 12'b111100000111;
            14'b01_001010111101: DATA = 12'b111100001000;
            14'b01_001010111110: DATA = 12'b111100001010;
            14'b01_001010111111: DATA = 12'b111100001011;
            14'b01_001011000000: DATA = 12'b111100001101;
            14'b01_001011000001: DATA = 12'b111100001110;
            14'b01_001011000010: DATA = 12'b111100010000;
            14'b01_001011000011: DATA = 12'b111100010001;
            14'b01_001011000100: DATA = 12'b111100010011;
            14'b01_001011000101: DATA = 12'b111100010100;
            14'b01_001011000110: DATA = 12'b111100010110;
            14'b01_001011000111: DATA = 12'b111100010111;
            14'b01_001011001000: DATA = 12'b111100011000;
            14'b01_001011001001: DATA = 12'b111100011010;
            14'b01_001011001010: DATA = 12'b111100011011;
            14'b01_001011001011: DATA = 12'b111100011101;
            14'b01_001011001100: DATA = 12'b111100011110;
            14'b01_001011001101: DATA = 12'b111100100000;
            14'b01_001011001110: DATA = 12'b111100100001;
            14'b01_001011001111: DATA = 12'b111100100011;
            14'b01_001011010000: DATA = 12'b111100100100;
            14'b01_001011010001: DATA = 12'b111100100101;
            14'b01_001011010010: DATA = 12'b111100100111;
            14'b01_001011010011: DATA = 12'b111100101000;
            14'b01_001011010100: DATA = 12'b111100101010;
            14'b01_001011010101: DATA = 12'b111100101011;
            14'b01_001011010110: DATA = 12'b111100101100;
            14'b01_001011010111: DATA = 12'b111100101110;
            14'b01_001011011000: DATA = 12'b111100101111;
            14'b01_001011011001: DATA = 12'b111100110000;
            14'b01_001011011010: DATA = 12'b111100110010;
            14'b01_001011011011: DATA = 12'b111100110011;
            14'b01_001011011100: DATA = 12'b111100110101;
            14'b01_001011011101: DATA = 12'b111100110110;
            14'b01_001011011110: DATA = 12'b111100110111;
            14'b01_001011011111: DATA = 12'b111100111001;
            14'b01_001011100000: DATA = 12'b111100111010;
            14'b01_001011100001: DATA = 12'b111100111011;
            14'b01_001011100010: DATA = 12'b111100111101;
            14'b01_001011100011: DATA = 12'b111100111110;
            14'b01_001011100100: DATA = 12'b111100111111;
            14'b01_001011100101: DATA = 12'b111101000001;
            14'b01_001011100110: DATA = 12'b111101000010;
            14'b01_001011100111: DATA = 12'b111101000011;
            14'b01_001011101000: DATA = 12'b111101000101;
            14'b01_001011101001: DATA = 12'b111101000110;
            14'b01_001011101010: DATA = 12'b111101000111;
            14'b01_001011101011: DATA = 12'b111101001000;
            14'b01_001011101100: DATA = 12'b111101001010;
            14'b01_001011101101: DATA = 12'b111101001011;
            14'b01_001011101110: DATA = 12'b111101001100;
            14'b01_001011101111: DATA = 12'b111101001110;
            14'b01_001011110000: DATA = 12'b111101001111;
            14'b01_001011110001: DATA = 12'b111101010000;
            14'b01_001011110010: DATA = 12'b111101010001;
            14'b01_001011110011: DATA = 12'b111101010011;
            14'b01_001011110100: DATA = 12'b111101010100;
            14'b01_001011110101: DATA = 12'b111101010101;
            14'b01_001011110110: DATA = 12'b111101010110;
            14'b01_001011110111: DATA = 12'b111101011000;
            14'b01_001011111000: DATA = 12'b111101011001;
            14'b01_001011111001: DATA = 12'b111101011010;
            14'b01_001011111010: DATA = 12'b111101011011;
            14'b01_001011111011: DATA = 12'b111101011101;
            14'b01_001011111100: DATA = 12'b111101011110;
            14'b01_001011111101: DATA = 12'b111101011111;
            14'b01_001011111110: DATA = 12'b111101100000;
            14'b01_001011111111: DATA = 12'b111101100001;
            14'b01_001100000000: DATA = 12'b111101100011;
            14'b01_001100000001: DATA = 12'b111101100100;
            14'b01_001100000010: DATA = 12'b111101100101;
            14'b01_001100000011: DATA = 12'b111101100110;
            14'b01_001100000100: DATA = 12'b111101100111;
            14'b01_001100000101: DATA = 12'b111101101001;
            14'b01_001100000110: DATA = 12'b111101101010;
            14'b01_001100000111: DATA = 12'b111101101011;
            14'b01_001100001000: DATA = 12'b111101101100;
            14'b01_001100001001: DATA = 12'b111101101101;
            14'b01_001100001010: DATA = 12'b111101101110;
            14'b01_001100001011: DATA = 12'b111101110000;
            14'b01_001100001100: DATA = 12'b111101110001;
            14'b01_001100001101: DATA = 12'b111101110010;
            14'b01_001100001110: DATA = 12'b111101110011;
            14'b01_001100001111: DATA = 12'b111101110100;
            14'b01_001100010000: DATA = 12'b111101110101;
            14'b01_001100010001: DATA = 12'b111101110110;
            14'b01_001100010010: DATA = 12'b111101111000;
            14'b01_001100010011: DATA = 12'b111101111001;
            14'b01_001100010100: DATA = 12'b111101111010;
            14'b01_001100010101: DATA = 12'b111101111011;
            14'b01_001100010110: DATA = 12'b111101111100;
            14'b01_001100010111: DATA = 12'b111101111101;
            14'b01_001100011000: DATA = 12'b111101111110;
            14'b01_001100011001: DATA = 12'b111101111111;
            14'b01_001100011010: DATA = 12'b111110000000;
            14'b01_001100011011: DATA = 12'b111110000001;
            14'b01_001100011100: DATA = 12'b111110000011;
            14'b01_001100011101: DATA = 12'b111110000100;
            14'b01_001100011110: DATA = 12'b111110000101;
            14'b01_001100011111: DATA = 12'b111110000110;
            14'b01_001100100000: DATA = 12'b111110000111;
            14'b01_001100100001: DATA = 12'b111110001000;
            14'b01_001100100010: DATA = 12'b111110001001;
            14'b01_001100100011: DATA = 12'b111110001010;
            14'b01_001100100100: DATA = 12'b111110001011;
            14'b01_001100100101: DATA = 12'b111110001100;
            14'b01_001100100110: DATA = 12'b111110001101;
            14'b01_001100100111: DATA = 12'b111110001110;
            14'b01_001100101000: DATA = 12'b111110001111;
            14'b01_001100101001: DATA = 12'b111110010000;
            14'b01_001100101010: DATA = 12'b111110010001;
            14'b01_001100101011: DATA = 12'b111110010010;
            14'b01_001100101100: DATA = 12'b111110010011;
            14'b01_001100101101: DATA = 12'b111110010100;
            14'b01_001100101110: DATA = 12'b111110010101;
            14'b01_001100101111: DATA = 12'b111110010110;
            14'b01_001100110000: DATA = 12'b111110010111;
            14'b01_001100110001: DATA = 12'b111110011000;
            14'b01_001100110010: DATA = 12'b111110011001;
            14'b01_001100110011: DATA = 12'b111110011010;
            14'b01_001100110100: DATA = 12'b111110011011;
            14'b01_001100110101: DATA = 12'b111110011100;
            14'b01_001100110110: DATA = 12'b111110011101;
            14'b01_001100110111: DATA = 12'b111110011110;
            14'b01_001100111000: DATA = 12'b111110011111;
            14'b01_001100111001: DATA = 12'b111110100000;
            14'b01_001100111010: DATA = 12'b111110100001;
            14'b01_001100111011: DATA = 12'b111110100010;
            14'b01_001100111100: DATA = 12'b111110100011;
            14'b01_001100111101: DATA = 12'b111110100100;
            14'b01_001100111110: DATA = 12'b111110100101;
            14'b01_001100111111: DATA = 12'b111110100101;
            14'b01_001101000000: DATA = 12'b111110100110;
            14'b01_001101000001: DATA = 12'b111110100111;
            14'b01_001101000010: DATA = 12'b111110101000;
            14'b01_001101000011: DATA = 12'b111110101001;
            14'b01_001101000100: DATA = 12'b111110101010;
            14'b01_001101000101: DATA = 12'b111110101011;
            14'b01_001101000110: DATA = 12'b111110101100;
            14'b01_001101000111: DATA = 12'b111110101101;
            14'b01_001101001000: DATA = 12'b111110101110;
            14'b01_001101001001: DATA = 12'b111110101110;
            14'b01_001101001010: DATA = 12'b111110101111;
            14'b01_001101001011: DATA = 12'b111110110000;
            14'b01_001101001100: DATA = 12'b111110110001;
            14'b01_001101001101: DATA = 12'b111110110010;
            14'b01_001101001110: DATA = 12'b111110110011;
            14'b01_001101001111: DATA = 12'b111110110100;
            14'b01_001101010000: DATA = 12'b111110110100;
            14'b01_001101010001: DATA = 12'b111110110101;
            14'b01_001101010010: DATA = 12'b111110110110;
            14'b01_001101010011: DATA = 12'b111110110111;
            14'b01_001101010100: DATA = 12'b111110111000;
            14'b01_001101010101: DATA = 12'b111110111000;
            14'b01_001101010110: DATA = 12'b111110111001;
            14'b01_001101010111: DATA = 12'b111110111010;
            14'b01_001101011000: DATA = 12'b111110111011;
            14'b01_001101011001: DATA = 12'b111110111100;
            14'b01_001101011010: DATA = 12'b111110111100;
            14'b01_001101011011: DATA = 12'b111110111101;
            14'b01_001101011100: DATA = 12'b111110111110;
            14'b01_001101011101: DATA = 12'b111110111111;
            14'b01_001101011110: DATA = 12'b111111000000;
            14'b01_001101011111: DATA = 12'b111111000000;
            14'b01_001101100000: DATA = 12'b111111000001;
            14'b01_001101100001: DATA = 12'b111111000010;
            14'b01_001101100010: DATA = 12'b111111000011;
            14'b01_001101100011: DATA = 12'b111111000011;
            14'b01_001101100100: DATA = 12'b111111000100;
            14'b01_001101100101: DATA = 12'b111111000101;
            14'b01_001101100110: DATA = 12'b111111000110;
            14'b01_001101100111: DATA = 12'b111111000110;
            14'b01_001101101000: DATA = 12'b111111000111;
            14'b01_001101101001: DATA = 12'b111111001000;
            14'b01_001101101010: DATA = 12'b111111001001;
            14'b01_001101101011: DATA = 12'b111111001001;
            14'b01_001101101100: DATA = 12'b111111001010;
            14'b01_001101101101: DATA = 12'b111111001011;
            14'b01_001101101110: DATA = 12'b111111001011;
            14'b01_001101101111: DATA = 12'b111111001100;
            14'b01_001101110000: DATA = 12'b111111001101;
            14'b01_001101110001: DATA = 12'b111111001101;
            14'b01_001101110010: DATA = 12'b111111001110;
            14'b01_001101110011: DATA = 12'b111111001111;
            14'b01_001101110100: DATA = 12'b111111001111;
            14'b01_001101110101: DATA = 12'b111111010000;
            14'b01_001101110110: DATA = 12'b111111010001;
            14'b01_001101110111: DATA = 12'b111111010001;
            14'b01_001101111000: DATA = 12'b111111010010;
            14'b01_001101111001: DATA = 12'b111111010011;
            14'b01_001101111010: DATA = 12'b111111010011;
            14'b01_001101111011: DATA = 12'b111111010100;
            14'b01_001101111100: DATA = 12'b111111010101;
            14'b01_001101111101: DATA = 12'b111111010101;
            14'b01_001101111110: DATA = 12'b111111010110;
            14'b01_001101111111: DATA = 12'b111111010111;
            14'b01_001110000000: DATA = 12'b111111010111;
            14'b01_001110000001: DATA = 12'b111111011000;
            14'b01_001110000010: DATA = 12'b111111011000;
            14'b01_001110000011: DATA = 12'b111111011001;
            14'b01_001110000100: DATA = 12'b111111011010;
            14'b01_001110000101: DATA = 12'b111111011010;
            14'b01_001110000110: DATA = 12'b111111011011;
            14'b01_001110000111: DATA = 12'b111111011011;
            14'b01_001110001000: DATA = 12'b111111011100;
            14'b01_001110001001: DATA = 12'b111111011100;
            14'b01_001110001010: DATA = 12'b111111011101;
            14'b01_001110001011: DATA = 12'b111111011110;
            14'b01_001110001100: DATA = 12'b111111011110;
            14'b01_001110001101: DATA = 12'b111111011111;
            14'b01_001110001110: DATA = 12'b111111011111;
            14'b01_001110001111: DATA = 12'b111111100000;
            14'b01_001110010000: DATA = 12'b111111100000;
            14'b01_001110010001: DATA = 12'b111111100001;
            14'b01_001110010010: DATA = 12'b111111100001;
            14'b01_001110010011: DATA = 12'b111111100010;
            14'b01_001110010100: DATA = 12'b111111100010;
            14'b01_001110010101: DATA = 12'b111111100011;
            14'b01_001110010110: DATA = 12'b111111100011;
            14'b01_001110010111: DATA = 12'b111111100100;
            14'b01_001110011000: DATA = 12'b111111100101;
            14'b01_001110011001: DATA = 12'b111111100101;
            14'b01_001110011010: DATA = 12'b111111100101;
            14'b01_001110011011: DATA = 12'b111111100110;
            14'b01_001110011100: DATA = 12'b111111100110;
            14'b01_001110011101: DATA = 12'b111111100111;
            14'b01_001110011110: DATA = 12'b111111100111;
            14'b01_001110011111: DATA = 12'b111111101000;
            14'b01_001110100000: DATA = 12'b111111101000;
            14'b01_001110100001: DATA = 12'b111111101001;
            14'b01_001110100010: DATA = 12'b111111101001;
            14'b01_001110100011: DATA = 12'b111111101010;
            14'b01_001110100100: DATA = 12'b111111101010;
            14'b01_001110100101: DATA = 12'b111111101011;
            14'b01_001110100110: DATA = 12'b111111101011;
            14'b01_001110100111: DATA = 12'b111111101011;
            14'b01_001110101000: DATA = 12'b111111101100;
            14'b01_001110101001: DATA = 12'b111111101100;
            14'b01_001110101010: DATA = 12'b111111101101;
            14'b01_001110101011: DATA = 12'b111111101101;
            14'b01_001110101100: DATA = 12'b111111101110;
            14'b01_001110101101: DATA = 12'b111111101110;
            14'b01_001110101110: DATA = 12'b111111101110;
            14'b01_001110101111: DATA = 12'b111111101111;
            14'b01_001110110000: DATA = 12'b111111101111;
            14'b01_001110110001: DATA = 12'b111111101111;
            14'b01_001110110010: DATA = 12'b111111110000;
            14'b01_001110110011: DATA = 12'b111111110000;
            14'b01_001110110100: DATA = 12'b111111110001;
            14'b01_001110110101: DATA = 12'b111111110001;
            14'b01_001110110110: DATA = 12'b111111110001;
            14'b01_001110110111: DATA = 12'b111111110010;
            14'b01_001110111000: DATA = 12'b111111110010;
            14'b01_001110111001: DATA = 12'b111111110010;
            14'b01_001110111010: DATA = 12'b111111110011;
            14'b01_001110111011: DATA = 12'b111111110011;
            14'b01_001110111100: DATA = 12'b111111110011;
            14'b01_001110111101: DATA = 12'b111111110100;
            14'b01_001110111110: DATA = 12'b111111110100;
            14'b01_001110111111: DATA = 12'b111111110100;
            14'b01_001111000000: DATA = 12'b111111110101;
            14'b01_001111000001: DATA = 12'b111111110101;
            14'b01_001111000010: DATA = 12'b111111110101;
            14'b01_001111000011: DATA = 12'b111111110110;
            14'b01_001111000100: DATA = 12'b111111110110;
            14'b01_001111000101: DATA = 12'b111111110110;
            14'b01_001111000110: DATA = 12'b111111110110;
            14'b01_001111000111: DATA = 12'b111111110111;
            14'b01_001111001000: DATA = 12'b111111110111;
            14'b01_001111001001: DATA = 12'b111111110111;
            14'b01_001111001010: DATA = 12'b111111110111;
            14'b01_001111001011: DATA = 12'b111111111000;
            14'b01_001111001100: DATA = 12'b111111111000;
            14'b01_001111001101: DATA = 12'b111111111000;
            14'b01_001111001110: DATA = 12'b111111111000;
            14'b01_001111001111: DATA = 12'b111111111001;
            14'b01_001111010000: DATA = 12'b111111111001;
            14'b01_001111010001: DATA = 12'b111111111001;
            14'b01_001111010010: DATA = 12'b111111111001;
            14'b01_001111010011: DATA = 12'b111111111010;
            14'b01_001111010100: DATA = 12'b111111111010;
            14'b01_001111010101: DATA = 12'b111111111010;
            14'b01_001111010110: DATA = 12'b111111111010;
            14'b01_001111010111: DATA = 12'b111111111010;
            14'b01_001111011000: DATA = 12'b111111111011;
            14'b01_001111011001: DATA = 12'b111111111011;
            14'b01_001111011010: DATA = 12'b111111111011;
            14'b01_001111011011: DATA = 12'b111111111011;
            14'b01_001111011100: DATA = 12'b111111111011;
            14'b01_001111011101: DATA = 12'b111111111100;
            14'b01_001111011110: DATA = 12'b111111111100;
            14'b01_001111011111: DATA = 12'b111111111100;
            14'b01_001111100000: DATA = 12'b111111111100;
            14'b01_001111100001: DATA = 12'b111111111100;
            14'b01_001111100010: DATA = 12'b111111111100;
            14'b01_001111100011: DATA = 12'b111111111100;
            14'b01_001111100100: DATA = 12'b111111111101;
            14'b01_001111100101: DATA = 12'b111111111101;
            14'b01_001111100110: DATA = 12'b111111111101;
            14'b01_001111100111: DATA = 12'b111111111101;
            14'b01_001111101000: DATA = 12'b111111111101;
            14'b01_001111101001: DATA = 12'b111111111101;
            14'b01_001111101010: DATA = 12'b111111111101;
            14'b01_001111101011: DATA = 12'b111111111101;
            14'b01_001111101100: DATA = 12'b111111111110;
            14'b01_001111101101: DATA = 12'b111111111110;
            14'b01_001111101110: DATA = 12'b111111111110;
            14'b01_001111101111: DATA = 12'b111111111110;
            14'b01_001111110000: DATA = 12'b111111111110;
            14'b01_001111110001: DATA = 12'b111111111110;
            14'b01_001111110010: DATA = 12'b111111111110;
            14'b01_001111110011: DATA = 12'b111111111110;
            14'b01_001111110100: DATA = 12'b111111111110;
            14'b01_001111110101: DATA = 12'b111111111110;
            14'b01_001111110110: DATA = 12'b111111111110;
            14'b01_001111110111: DATA = 12'b111111111110;
            14'b01_001111111000: DATA = 12'b111111111110;
            14'b01_001111111001: DATA = 12'b111111111110;
            14'b01_001111111010: DATA = 12'b111111111110;
            14'b01_001111111011: DATA = 12'b111111111110;
            14'b01_001111111100: DATA = 12'b111111111110;
            14'b01_001111111101: DATA = 12'b111111111110;
            14'b01_001111111110: DATA = 12'b111111111110;
            14'b01_001111111111: DATA = 12'b111111111110;
            14'b01_010000000000: DATA = 12'b111111111111;
            14'b01_010000000001: DATA = 12'b111111111110;
            14'b01_010000000010: DATA = 12'b111111111110;
            14'b01_010000000011: DATA = 12'b111111111110;
            14'b01_010000000100: DATA = 12'b111111111110;
            14'b01_010000000101: DATA = 12'b111111111110;
            14'b01_010000000110: DATA = 12'b111111111110;
            14'b01_010000000111: DATA = 12'b111111111110;
            14'b01_010000001000: DATA = 12'b111111111110;
            14'b01_010000001001: DATA = 12'b111111111110;
            14'b01_010000001010: DATA = 12'b111111111110;
            14'b01_010000001011: DATA = 12'b111111111110;
            14'b01_010000001100: DATA = 12'b111111111110;
            14'b01_010000001101: DATA = 12'b111111111110;
            14'b01_010000001110: DATA = 12'b111111111110;
            14'b01_010000001111: DATA = 12'b111111111110;
            14'b01_010000010000: DATA = 12'b111111111110;
            14'b01_010000010001: DATA = 12'b111111111110;
            14'b01_010000010010: DATA = 12'b111111111110;
            14'b01_010000010011: DATA = 12'b111111111110;
            14'b01_010000010100: DATA = 12'b111111111110;
            14'b01_010000010101: DATA = 12'b111111111101;
            14'b01_010000010110: DATA = 12'b111111111101;
            14'b01_010000010111: DATA = 12'b111111111101;
            14'b01_010000011000: DATA = 12'b111111111101;
            14'b01_010000011001: DATA = 12'b111111111101;
            14'b01_010000011010: DATA = 12'b111111111101;
            14'b01_010000011011: DATA = 12'b111111111101;
            14'b01_010000011100: DATA = 12'b111111111101;
            14'b01_010000011101: DATA = 12'b111111111100;
            14'b01_010000011110: DATA = 12'b111111111100;
            14'b01_010000011111: DATA = 12'b111111111100;
            14'b01_010000100000: DATA = 12'b111111111100;
            14'b01_010000100001: DATA = 12'b111111111100;
            14'b01_010000100010: DATA = 12'b111111111100;
            14'b01_010000100011: DATA = 12'b111111111100;
            14'b01_010000100100: DATA = 12'b111111111011;
            14'b01_010000100101: DATA = 12'b111111111011;
            14'b01_010000100110: DATA = 12'b111111111011;
            14'b01_010000100111: DATA = 12'b111111111011;
            14'b01_010000101000: DATA = 12'b111111111011;
            14'b01_010000101001: DATA = 12'b111111111010;
            14'b01_010000101010: DATA = 12'b111111111010;
            14'b01_010000101011: DATA = 12'b111111111010;
            14'b01_010000101100: DATA = 12'b111111111010;
            14'b01_010000101101: DATA = 12'b111111111010;
            14'b01_010000101110: DATA = 12'b111111111001;
            14'b01_010000101111: DATA = 12'b111111111001;
            14'b01_010000110000: DATA = 12'b111111111001;
            14'b01_010000110001: DATA = 12'b111111111001;
            14'b01_010000110010: DATA = 12'b111111111000;
            14'b01_010000110011: DATA = 12'b111111111000;
            14'b01_010000110100: DATA = 12'b111111111000;
            14'b01_010000110101: DATA = 12'b111111111000;
            14'b01_010000110110: DATA = 12'b111111110111;
            14'b01_010000110111: DATA = 12'b111111110111;
            14'b01_010000111000: DATA = 12'b111111110111;
            14'b01_010000111001: DATA = 12'b111111110111;
            14'b01_010000111010: DATA = 12'b111111110110;
            14'b01_010000111011: DATA = 12'b111111110110;
            14'b01_010000111100: DATA = 12'b111111110110;
            14'b01_010000111101: DATA = 12'b111111110110;
            14'b01_010000111110: DATA = 12'b111111110101;
            14'b01_010000111111: DATA = 12'b111111110101;
            14'b01_010001000000: DATA = 12'b111111110101;
            14'b01_010001000001: DATA = 12'b111111110100;
            14'b01_010001000010: DATA = 12'b111111110100;
            14'b01_010001000011: DATA = 12'b111111110100;
            14'b01_010001000100: DATA = 12'b111111110011;
            14'b01_010001000101: DATA = 12'b111111110011;
            14'b01_010001000110: DATA = 12'b111111110011;
            14'b01_010001000111: DATA = 12'b111111110010;
            14'b01_010001001000: DATA = 12'b111111110010;
            14'b01_010001001001: DATA = 12'b111111110010;
            14'b01_010001001010: DATA = 12'b111111110001;
            14'b01_010001001011: DATA = 12'b111111110001;
            14'b01_010001001100: DATA = 12'b111111110001;
            14'b01_010001001101: DATA = 12'b111111110000;
            14'b01_010001001110: DATA = 12'b111111110000;
            14'b01_010001001111: DATA = 12'b111111101111;
            14'b01_010001010000: DATA = 12'b111111101111;
            14'b01_010001010001: DATA = 12'b111111101111;
            14'b01_010001010010: DATA = 12'b111111101110;
            14'b01_010001010011: DATA = 12'b111111101110;
            14'b01_010001010100: DATA = 12'b111111101110;
            14'b01_010001010101: DATA = 12'b111111101101;
            14'b01_010001010110: DATA = 12'b111111101101;
            14'b01_010001010111: DATA = 12'b111111101100;
            14'b01_010001011000: DATA = 12'b111111101100;
            14'b01_010001011001: DATA = 12'b111111101011;
            14'b01_010001011010: DATA = 12'b111111101011;
            14'b01_010001011011: DATA = 12'b111111101011;
            14'b01_010001011100: DATA = 12'b111111101010;
            14'b01_010001011101: DATA = 12'b111111101010;
            14'b01_010001011110: DATA = 12'b111111101001;
            14'b01_010001011111: DATA = 12'b111111101001;
            14'b01_010001100000: DATA = 12'b111111101000;
            14'b01_010001100001: DATA = 12'b111111101000;
            14'b01_010001100010: DATA = 12'b111111100111;
            14'b01_010001100011: DATA = 12'b111111100111;
            14'b01_010001100100: DATA = 12'b111111100110;
            14'b01_010001100101: DATA = 12'b111111100110;
            14'b01_010001100110: DATA = 12'b111111100101;
            14'b01_010001100111: DATA = 12'b111111100101;
            14'b01_010001101000: DATA = 12'b111111100101;
            14'b01_010001101001: DATA = 12'b111111100100;
            14'b01_010001101010: DATA = 12'b111111100011;
            14'b01_010001101011: DATA = 12'b111111100011;
            14'b01_010001101100: DATA = 12'b111111100010;
            14'b01_010001101101: DATA = 12'b111111100010;
            14'b01_010001101110: DATA = 12'b111111100001;
            14'b01_010001101111: DATA = 12'b111111100001;
            14'b01_010001110000: DATA = 12'b111111100000;
            14'b01_010001110001: DATA = 12'b111111100000;
            14'b01_010001110010: DATA = 12'b111111011111;
            14'b01_010001110011: DATA = 12'b111111011111;
            14'b01_010001110100: DATA = 12'b111111011110;
            14'b01_010001110101: DATA = 12'b111111011110;
            14'b01_010001110110: DATA = 12'b111111011101;
            14'b01_010001110111: DATA = 12'b111111011100;
            14'b01_010001111000: DATA = 12'b111111011100;
            14'b01_010001111001: DATA = 12'b111111011011;
            14'b01_010001111010: DATA = 12'b111111011011;
            14'b01_010001111011: DATA = 12'b111111011010;
            14'b01_010001111100: DATA = 12'b111111011010;
            14'b01_010001111101: DATA = 12'b111111011001;
            14'b01_010001111110: DATA = 12'b111111011000;
            14'b01_010001111111: DATA = 12'b111111011000;
            14'b01_010010000000: DATA = 12'b111111010111;
            14'b01_010010000001: DATA = 12'b111111010111;
            14'b01_010010000010: DATA = 12'b111111010110;
            14'b01_010010000011: DATA = 12'b111111010101;
            14'b01_010010000100: DATA = 12'b111111010101;
            14'b01_010010000101: DATA = 12'b111111010100;
            14'b01_010010000110: DATA = 12'b111111010011;
            14'b01_010010000111: DATA = 12'b111111010011;
            14'b01_010010001000: DATA = 12'b111111010010;
            14'b01_010010001001: DATA = 12'b111111010001;
            14'b01_010010001010: DATA = 12'b111111010001;
            14'b01_010010001011: DATA = 12'b111111010000;
            14'b01_010010001100: DATA = 12'b111111001111;
            14'b01_010010001101: DATA = 12'b111111001111;
            14'b01_010010001110: DATA = 12'b111111001110;
            14'b01_010010001111: DATA = 12'b111111001101;
            14'b01_010010010000: DATA = 12'b111111001101;
            14'b01_010010010001: DATA = 12'b111111001100;
            14'b01_010010010010: DATA = 12'b111111001011;
            14'b01_010010010011: DATA = 12'b111111001011;
            14'b01_010010010100: DATA = 12'b111111001010;
            14'b01_010010010101: DATA = 12'b111111001001;
            14'b01_010010010110: DATA = 12'b111111001001;
            14'b01_010010010111: DATA = 12'b111111001000;
            14'b01_010010011000: DATA = 12'b111111000111;
            14'b01_010010011001: DATA = 12'b111111000110;
            14'b01_010010011010: DATA = 12'b111111000110;
            14'b01_010010011011: DATA = 12'b111111000101;
            14'b01_010010011100: DATA = 12'b111111000100;
            14'b01_010010011101: DATA = 12'b111111000011;
            14'b01_010010011110: DATA = 12'b111111000011;
            14'b01_010010011111: DATA = 12'b111111000010;
            14'b01_010010100000: DATA = 12'b111111000001;
            14'b01_010010100001: DATA = 12'b111111000000;
            14'b01_010010100010: DATA = 12'b111111000000;
            14'b01_010010100011: DATA = 12'b111110111111;
            14'b01_010010100100: DATA = 12'b111110111110;
            14'b01_010010100101: DATA = 12'b111110111101;
            14'b01_010010100110: DATA = 12'b111110111100;
            14'b01_010010100111: DATA = 12'b111110111100;
            14'b01_010010101000: DATA = 12'b111110111011;
            14'b01_010010101001: DATA = 12'b111110111010;
            14'b01_010010101010: DATA = 12'b111110111001;
            14'b01_010010101011: DATA = 12'b111110111000;
            14'b01_010010101100: DATA = 12'b111110111000;
            14'b01_010010101101: DATA = 12'b111110110111;
            14'b01_010010101110: DATA = 12'b111110110110;
            14'b01_010010101111: DATA = 12'b111110110101;
            14'b01_010010110000: DATA = 12'b111110110100;
            14'b01_010010110001: DATA = 12'b111110110100;
            14'b01_010010110010: DATA = 12'b111110110011;
            14'b01_010010110011: DATA = 12'b111110110010;
            14'b01_010010110100: DATA = 12'b111110110001;
            14'b01_010010110101: DATA = 12'b111110110000;
            14'b01_010010110110: DATA = 12'b111110101111;
            14'b01_010010110111: DATA = 12'b111110101110;
            14'b01_010010111000: DATA = 12'b111110101110;
            14'b01_010010111001: DATA = 12'b111110101101;
            14'b01_010010111010: DATA = 12'b111110101100;
            14'b01_010010111011: DATA = 12'b111110101011;
            14'b01_010010111100: DATA = 12'b111110101010;
            14'b01_010010111101: DATA = 12'b111110101001;
            14'b01_010010111110: DATA = 12'b111110101000;
            14'b01_010010111111: DATA = 12'b111110100111;
            14'b01_010011000000: DATA = 12'b111110100110;
            14'b01_010011000001: DATA = 12'b111110100101;
            14'b01_010011000010: DATA = 12'b111110100101;
            14'b01_010011000011: DATA = 12'b111110100100;
            14'b01_010011000100: DATA = 12'b111110100011;
            14'b01_010011000101: DATA = 12'b111110100010;
            14'b01_010011000110: DATA = 12'b111110100001;
            14'b01_010011000111: DATA = 12'b111110100000;
            14'b01_010011001000: DATA = 12'b111110011111;
            14'b01_010011001001: DATA = 12'b111110011110;
            14'b01_010011001010: DATA = 12'b111110011101;
            14'b01_010011001011: DATA = 12'b111110011100;
            14'b01_010011001100: DATA = 12'b111110011011;
            14'b01_010011001101: DATA = 12'b111110011010;
            14'b01_010011001110: DATA = 12'b111110011001;
            14'b01_010011001111: DATA = 12'b111110011000;
            14'b01_010011010000: DATA = 12'b111110010111;
            14'b01_010011010001: DATA = 12'b111110010110;
            14'b01_010011010010: DATA = 12'b111110010101;
            14'b01_010011010011: DATA = 12'b111110010100;
            14'b01_010011010100: DATA = 12'b111110010011;
            14'b01_010011010101: DATA = 12'b111110010010;
            14'b01_010011010110: DATA = 12'b111110010001;
            14'b01_010011010111: DATA = 12'b111110010000;
            14'b01_010011011000: DATA = 12'b111110001111;
            14'b01_010011011001: DATA = 12'b111110001110;
            14'b01_010011011010: DATA = 12'b111110001101;
            14'b01_010011011011: DATA = 12'b111110001100;
            14'b01_010011011100: DATA = 12'b111110001011;
            14'b01_010011011101: DATA = 12'b111110001010;
            14'b01_010011011110: DATA = 12'b111110001001;
            14'b01_010011011111: DATA = 12'b111110001000;
            14'b01_010011100000: DATA = 12'b111110000111;
            14'b01_010011100001: DATA = 12'b111110000110;
            14'b01_010011100010: DATA = 12'b111110000101;
            14'b01_010011100011: DATA = 12'b111110000100;
            14'b01_010011100100: DATA = 12'b111110000011;
            14'b01_010011100101: DATA = 12'b111110000001;
            14'b01_010011100110: DATA = 12'b111110000000;
            14'b01_010011100111: DATA = 12'b111101111111;
            14'b01_010011101000: DATA = 12'b111101111110;
            14'b01_010011101001: DATA = 12'b111101111101;
            14'b01_010011101010: DATA = 12'b111101111100;
            14'b01_010011101011: DATA = 12'b111101111011;
            14'b01_010011101100: DATA = 12'b111101111010;
            14'b01_010011101101: DATA = 12'b111101111001;
            14'b01_010011101110: DATA = 12'b111101111000;
            14'b01_010011101111: DATA = 12'b111101110110;
            14'b01_010011110000: DATA = 12'b111101110101;
            14'b01_010011110001: DATA = 12'b111101110100;
            14'b01_010011110010: DATA = 12'b111101110011;
            14'b01_010011110011: DATA = 12'b111101110010;
            14'b01_010011110100: DATA = 12'b111101110001;
            14'b01_010011110101: DATA = 12'b111101110000;
            14'b01_010011110110: DATA = 12'b111101101110;
            14'b01_010011110111: DATA = 12'b111101101101;
            14'b01_010011111000: DATA = 12'b111101101100;
            14'b01_010011111001: DATA = 12'b111101101011;
            14'b01_010011111010: DATA = 12'b111101101010;
            14'b01_010011111011: DATA = 12'b111101101001;
            14'b01_010011111100: DATA = 12'b111101100111;
            14'b01_010011111101: DATA = 12'b111101100110;
            14'b01_010011111110: DATA = 12'b111101100101;
            14'b01_010011111111: DATA = 12'b111101100100;
            14'b01_010100000000: DATA = 12'b111101100011;
            14'b01_010100000001: DATA = 12'b111101100001;
            14'b01_010100000010: DATA = 12'b111101100000;
            14'b01_010100000011: DATA = 12'b111101011111;
            14'b01_010100000100: DATA = 12'b111101011110;
            14'b01_010100000101: DATA = 12'b111101011101;
            14'b01_010100000110: DATA = 12'b111101011011;
            14'b01_010100000111: DATA = 12'b111101011010;
            14'b01_010100001000: DATA = 12'b111101011001;
            14'b01_010100001001: DATA = 12'b111101011000;
            14'b01_010100001010: DATA = 12'b111101010110;
            14'b01_010100001011: DATA = 12'b111101010101;
            14'b01_010100001100: DATA = 12'b111101010100;
            14'b01_010100001101: DATA = 12'b111101010011;
            14'b01_010100001110: DATA = 12'b111101010001;
            14'b01_010100001111: DATA = 12'b111101010000;
            14'b01_010100010000: DATA = 12'b111101001111;
            14'b01_010100010001: DATA = 12'b111101001110;
            14'b01_010100010010: DATA = 12'b111101001100;
            14'b01_010100010011: DATA = 12'b111101001011;
            14'b01_010100010100: DATA = 12'b111101001010;
            14'b01_010100010101: DATA = 12'b111101001000;
            14'b01_010100010110: DATA = 12'b111101000111;
            14'b01_010100010111: DATA = 12'b111101000110;
            14'b01_010100011000: DATA = 12'b111101000101;
            14'b01_010100011001: DATA = 12'b111101000011;
            14'b01_010100011010: DATA = 12'b111101000010;
            14'b01_010100011011: DATA = 12'b111101000001;
            14'b01_010100011100: DATA = 12'b111100111111;
            14'b01_010100011101: DATA = 12'b111100111110;
            14'b01_010100011110: DATA = 12'b111100111101;
            14'b01_010100011111: DATA = 12'b111100111011;
            14'b01_010100100000: DATA = 12'b111100111010;
            14'b01_010100100001: DATA = 12'b111100111001;
            14'b01_010100100010: DATA = 12'b111100110111;
            14'b01_010100100011: DATA = 12'b111100110110;
            14'b01_010100100100: DATA = 12'b111100110101;
            14'b01_010100100101: DATA = 12'b111100110011;
            14'b01_010100100110: DATA = 12'b111100110010;
            14'b01_010100100111: DATA = 12'b111100110000;
            14'b01_010100101000: DATA = 12'b111100101111;
            14'b01_010100101001: DATA = 12'b111100101110;
            14'b01_010100101010: DATA = 12'b111100101100;
            14'b01_010100101011: DATA = 12'b111100101011;
            14'b01_010100101100: DATA = 12'b111100101010;
            14'b01_010100101101: DATA = 12'b111100101000;
            14'b01_010100101110: DATA = 12'b111100100111;
            14'b01_010100101111: DATA = 12'b111100100101;
            14'b01_010100110000: DATA = 12'b111100100100;
            14'b01_010100110001: DATA = 12'b111100100011;
            14'b01_010100110010: DATA = 12'b111100100001;
            14'b01_010100110011: DATA = 12'b111100100000;
            14'b01_010100110100: DATA = 12'b111100011110;
            14'b01_010100110101: DATA = 12'b111100011101;
            14'b01_010100110110: DATA = 12'b111100011011;
            14'b01_010100110111: DATA = 12'b111100011010;
            14'b01_010100111000: DATA = 12'b111100011000;
            14'b01_010100111001: DATA = 12'b111100010111;
            14'b01_010100111010: DATA = 12'b111100010110;
            14'b01_010100111011: DATA = 12'b111100010100;
            14'b01_010100111100: DATA = 12'b111100010011;
            14'b01_010100111101: DATA = 12'b111100010001;
            14'b01_010100111110: DATA = 12'b111100010000;
            14'b01_010100111111: DATA = 12'b111100001110;
            14'b01_010101000000: DATA = 12'b111100001101;
            14'b01_010101000001: DATA = 12'b111100001011;
            14'b01_010101000010: DATA = 12'b111100001010;
            14'b01_010101000011: DATA = 12'b111100001000;
            14'b01_010101000100: DATA = 12'b111100000111;
            14'b01_010101000101: DATA = 12'b111100000101;
            14'b01_010101000110: DATA = 12'b111100000100;
            14'b01_010101000111: DATA = 12'b111100000010;
            14'b01_010101001000: DATA = 12'b111100000001;
            14'b01_010101001001: DATA = 12'b111011111111;
            14'b01_010101001010: DATA = 12'b111011111110;
            14'b01_010101001011: DATA = 12'b111011111100;
            14'b01_010101001100: DATA = 12'b111011111011;
            14'b01_010101001101: DATA = 12'b111011111001;
            14'b01_010101001110: DATA = 12'b111011111000;
            14'b01_010101001111: DATA = 12'b111011110110;
            14'b01_010101010000: DATA = 12'b111011110101;
            14'b01_010101010001: DATA = 12'b111011110011;
            14'b01_010101010010: DATA = 12'b111011110001;
            14'b01_010101010011: DATA = 12'b111011110000;
            14'b01_010101010100: DATA = 12'b111011101110;
            14'b01_010101010101: DATA = 12'b111011101101;
            14'b01_010101010110: DATA = 12'b111011101011;
            14'b01_010101010111: DATA = 12'b111011101010;
            14'b01_010101011000: DATA = 12'b111011101000;
            14'b01_010101011001: DATA = 12'b111011100110;
            14'b01_010101011010: DATA = 12'b111011100101;
            14'b01_010101011011: DATA = 12'b111011100011;
            14'b01_010101011100: DATA = 12'b111011100010;
            14'b01_010101011101: DATA = 12'b111011100000;
            14'b01_010101011110: DATA = 12'b111011011110;
            14'b01_010101011111: DATA = 12'b111011011101;
            14'b01_010101100000: DATA = 12'b111011011011;
            14'b01_010101100001: DATA = 12'b111011011010;
            14'b01_010101100010: DATA = 12'b111011011000;
            14'b01_010101100011: DATA = 12'b111011010110;
            14'b01_010101100100: DATA = 12'b111011010101;
            14'b01_010101100101: DATA = 12'b111011010011;
            14'b01_010101100110: DATA = 12'b111011010010;
            14'b01_010101100111: DATA = 12'b111011010000;
            14'b01_010101101000: DATA = 12'b111011001110;
            14'b01_010101101001: DATA = 12'b111011001101;
            14'b01_010101101010: DATA = 12'b111011001011;
            14'b01_010101101011: DATA = 12'b111011001001;
            14'b01_010101101100: DATA = 12'b111011001000;
            14'b01_010101101101: DATA = 12'b111011000110;
            14'b01_010101101110: DATA = 12'b111011000100;
            14'b01_010101101111: DATA = 12'b111011000011;
            14'b01_010101110000: DATA = 12'b111011000001;
            14'b01_010101110001: DATA = 12'b111010111111;
            14'b01_010101110010: DATA = 12'b111010111110;
            14'b01_010101110011: DATA = 12'b111010111100;
            14'b01_010101110100: DATA = 12'b111010111010;
            14'b01_010101110101: DATA = 12'b111010111000;
            14'b01_010101110110: DATA = 12'b111010110111;
            14'b01_010101110111: DATA = 12'b111010110101;
            14'b01_010101111000: DATA = 12'b111010110011;
            14'b01_010101111001: DATA = 12'b111010110010;
            14'b01_010101111010: DATA = 12'b111010110000;
            14'b01_010101111011: DATA = 12'b111010101110;
            14'b01_010101111100: DATA = 12'b111010101100;
            14'b01_010101111101: DATA = 12'b111010101011;
            14'b01_010101111110: DATA = 12'b111010101001;
            14'b01_010101111111: DATA = 12'b111010100111;
            14'b01_010110000000: DATA = 12'b111010100110;
            14'b01_010110000001: DATA = 12'b111010100100;
            14'b01_010110000010: DATA = 12'b111010100010;
            14'b01_010110000011: DATA = 12'b111010100000;
            14'b01_010110000100: DATA = 12'b111010011111;
            14'b01_010110000101: DATA = 12'b111010011101;
            14'b01_010110000110: DATA = 12'b111010011011;
            14'b01_010110000111: DATA = 12'b111010011001;
            14'b01_010110001000: DATA = 12'b111010010111;
            14'b01_010110001001: DATA = 12'b111010010110;
            14'b01_010110001010: DATA = 12'b111010010100;
            14'b01_010110001011: DATA = 12'b111010010010;
            14'b01_010110001100: DATA = 12'b111010010000;
            14'b01_010110001101: DATA = 12'b111010001111;
            14'b01_010110001110: DATA = 12'b111010001101;
            14'b01_010110001111: DATA = 12'b111010001011;
            14'b01_010110010000: DATA = 12'b111010001001;
            14'b01_010110010001: DATA = 12'b111010000111;
            14'b01_010110010010: DATA = 12'b111010000101;
            14'b01_010110010011: DATA = 12'b111010000100;
            14'b01_010110010100: DATA = 12'b111010000010;
            14'b01_010110010101: DATA = 12'b111010000000;
            14'b01_010110010110: DATA = 12'b111001111110;
            14'b01_010110010111: DATA = 12'b111001111100;
            14'b01_010110011000: DATA = 12'b111001111011;
            14'b01_010110011001: DATA = 12'b111001111001;
            14'b01_010110011010: DATA = 12'b111001110111;
            14'b01_010110011011: DATA = 12'b111001110101;
            14'b01_010110011100: DATA = 12'b111001110011;
            14'b01_010110011101: DATA = 12'b111001110001;
            14'b01_010110011110: DATA = 12'b111001101111;
            14'b01_010110011111: DATA = 12'b111001101110;
            14'b01_010110100000: DATA = 12'b111001101100;
            14'b01_010110100001: DATA = 12'b111001101010;
            14'b01_010110100010: DATA = 12'b111001101000;
            14'b01_010110100011: DATA = 12'b111001100110;
            14'b01_010110100100: DATA = 12'b111001100100;
            14'b01_010110100101: DATA = 12'b111001100010;
            14'b01_010110100110: DATA = 12'b111001100000;
            14'b01_010110100111: DATA = 12'b111001011110;
            14'b01_010110101000: DATA = 12'b111001011101;
            14'b01_010110101001: DATA = 12'b111001011011;
            14'b01_010110101010: DATA = 12'b111001011001;
            14'b01_010110101011: DATA = 12'b111001010111;
            14'b01_010110101100: DATA = 12'b111001010101;
            14'b01_010110101101: DATA = 12'b111001010011;
            14'b01_010110101110: DATA = 12'b111001010001;
            14'b01_010110101111: DATA = 12'b111001001111;
            14'b01_010110110000: DATA = 12'b111001001101;
            14'b01_010110110001: DATA = 12'b111001001011;
            14'b01_010110110010: DATA = 12'b111001001001;
            14'b01_010110110011: DATA = 12'b111001000111;
            14'b01_010110110100: DATA = 12'b111001000101;
            14'b01_010110110101: DATA = 12'b111001000100;
            14'b01_010110110110: DATA = 12'b111001000010;
            14'b01_010110110111: DATA = 12'b111001000000;
            14'b01_010110111000: DATA = 12'b111000111110;
            14'b01_010110111001: DATA = 12'b111000111100;
            14'b01_010110111010: DATA = 12'b111000111010;
            14'b01_010110111011: DATA = 12'b111000111000;
            14'b01_010110111100: DATA = 12'b111000110110;
            14'b01_010110111101: DATA = 12'b111000110100;
            14'b01_010110111110: DATA = 12'b111000110010;
            14'b01_010110111111: DATA = 12'b111000110000;
            14'b01_010111000000: DATA = 12'b111000101110;
            14'b01_010111000001: DATA = 12'b111000101100;
            14'b01_010111000010: DATA = 12'b111000101010;
            14'b01_010111000011: DATA = 12'b111000101000;
            14'b01_010111000100: DATA = 12'b111000100110;
            14'b01_010111000101: DATA = 12'b111000100100;
            14'b01_010111000110: DATA = 12'b111000100010;
            14'b01_010111000111: DATA = 12'b111000100000;
            14'b01_010111001000: DATA = 12'b111000011110;
            14'b01_010111001001: DATA = 12'b111000011100;
            14'b01_010111001010: DATA = 12'b111000011010;
            14'b01_010111001011: DATA = 12'b111000011000;
            14'b01_010111001100: DATA = 12'b111000010110;
            14'b01_010111001101: DATA = 12'b111000010100;
            14'b01_010111001110: DATA = 12'b111000010010;
            14'b01_010111001111: DATA = 12'b111000010000;
            14'b01_010111010000: DATA = 12'b111000001110;
            14'b01_010111010001: DATA = 12'b111000001011;
            14'b01_010111010010: DATA = 12'b111000001001;
            14'b01_010111010011: DATA = 12'b111000000111;
            14'b01_010111010100: DATA = 12'b111000000101;
            14'b01_010111010101: DATA = 12'b111000000011;
            14'b01_010111010110: DATA = 12'b111000000001;
            14'b01_010111010111: DATA = 12'b110111111111;
            14'b01_010111011000: DATA = 12'b110111111101;
            14'b01_010111011001: DATA = 12'b110111111011;
            14'b01_010111011010: DATA = 12'b110111111001;
            14'b01_010111011011: DATA = 12'b110111110111;
            14'b01_010111011100: DATA = 12'b110111110101;
            14'b01_010111011101: DATA = 12'b110111110011;
            14'b01_010111011110: DATA = 12'b110111110000;
            14'b01_010111011111: DATA = 12'b110111101110;
            14'b01_010111100000: DATA = 12'b110111101100;
            14'b01_010111100001: DATA = 12'b110111101010;
            14'b01_010111100010: DATA = 12'b110111101000;
            14'b01_010111100011: DATA = 12'b110111100110;
            14'b01_010111100100: DATA = 12'b110111100100;
            14'b01_010111100101: DATA = 12'b110111100010;
            14'b01_010111100110: DATA = 12'b110111100000;
            14'b01_010111100111: DATA = 12'b110111011101;
            14'b01_010111101000: DATA = 12'b110111011011;
            14'b01_010111101001: DATA = 12'b110111011001;
            14'b01_010111101010: DATA = 12'b110111010111;
            14'b01_010111101011: DATA = 12'b110111010101;
            14'b01_010111101100: DATA = 12'b110111010011;
            14'b01_010111101101: DATA = 12'b110111010001;
            14'b01_010111101110: DATA = 12'b110111001110;
            14'b01_010111101111: DATA = 12'b110111001100;
            14'b01_010111110000: DATA = 12'b110111001010;
            14'b01_010111110001: DATA = 12'b110111001000;
            14'b01_010111110010: DATA = 12'b110111000110;
            14'b01_010111110011: DATA = 12'b110111000100;
            14'b01_010111110100: DATA = 12'b110111000001;
            14'b01_010111110101: DATA = 12'b110110111111;
            14'b01_010111110110: DATA = 12'b110110111101;
            14'b01_010111110111: DATA = 12'b110110111011;
            14'b01_010111111000: DATA = 12'b110110111001;
            14'b01_010111111001: DATA = 12'b110110110110;
            14'b01_010111111010: DATA = 12'b110110110100;
            14'b01_010111111011: DATA = 12'b110110110010;
            14'b01_010111111100: DATA = 12'b110110110000;
            14'b01_010111111101: DATA = 12'b110110101110;
            14'b01_010111111110: DATA = 12'b110110101011;
            14'b01_010111111111: DATA = 12'b110110101001;
            14'b01_011000000000: DATA = 12'b110110100111;
            14'b01_011000000001: DATA = 12'b110110100101;
            14'b01_011000000010: DATA = 12'b110110100011;
            14'b01_011000000011: DATA = 12'b110110100000;
            14'b01_011000000100: DATA = 12'b110110011110;
            14'b01_011000000101: DATA = 12'b110110011100;
            14'b01_011000000110: DATA = 12'b110110011010;
            14'b01_011000000111: DATA = 12'b110110010111;
            14'b01_011000001000: DATA = 12'b110110010101;
            14'b01_011000001001: DATA = 12'b110110010011;
            14'b01_011000001010: DATA = 12'b110110010001;
            14'b01_011000001011: DATA = 12'b110110001110;
            14'b01_011000001100: DATA = 12'b110110001100;
            14'b01_011000001101: DATA = 12'b110110001010;
            14'b01_011000001110: DATA = 12'b110110001000;
            14'b01_011000001111: DATA = 12'b110110000101;
            14'b01_011000010000: DATA = 12'b110110000011;
            14'b01_011000010001: DATA = 12'b110110000001;
            14'b01_011000010010: DATA = 12'b110101111110;
            14'b01_011000010011: DATA = 12'b110101111100;
            14'b01_011000010100: DATA = 12'b110101111010;
            14'b01_011000010101: DATA = 12'b110101111000;
            14'b01_011000010110: DATA = 12'b110101110101;
            14'b01_011000010111: DATA = 12'b110101110011;
            14'b01_011000011000: DATA = 12'b110101110001;
            14'b01_011000011001: DATA = 12'b110101101110;
            14'b01_011000011010: DATA = 12'b110101101100;
            14'b01_011000011011: DATA = 12'b110101101010;
            14'b01_011000011100: DATA = 12'b110101100111;
            14'b01_011000011101: DATA = 12'b110101100101;
            14'b01_011000011110: DATA = 12'b110101100011;
            14'b01_011000011111: DATA = 12'b110101100001;
            14'b01_011000100000: DATA = 12'b110101011110;
            14'b01_011000100001: DATA = 12'b110101011100;
            14'b01_011000100010: DATA = 12'b110101011010;
            14'b01_011000100011: DATA = 12'b110101010111;
            14'b01_011000100100: DATA = 12'b110101010101;
            14'b01_011000100101: DATA = 12'b110101010011;
            14'b01_011000100110: DATA = 12'b110101010000;
            14'b01_011000100111: DATA = 12'b110101001110;
            14'b01_011000101000: DATA = 12'b110101001011;
            14'b01_011000101001: DATA = 12'b110101001001;
            14'b01_011000101010: DATA = 12'b110101000111;
            14'b01_011000101011: DATA = 12'b110101000100;
            14'b01_011000101100: DATA = 12'b110101000010;
            14'b01_011000101101: DATA = 12'b110101000000;
            14'b01_011000101110: DATA = 12'b110100111101;
            14'b01_011000101111: DATA = 12'b110100111011;
            14'b01_011000110000: DATA = 12'b110100111001;
            14'b01_011000110001: DATA = 12'b110100110110;
            14'b01_011000110010: DATA = 12'b110100110100;
            14'b01_011000110011: DATA = 12'b110100110001;
            14'b01_011000110100: DATA = 12'b110100101111;
            14'b01_011000110101: DATA = 12'b110100101101;
            14'b01_011000110110: DATA = 12'b110100101010;
            14'b01_011000110111: DATA = 12'b110100101000;
            14'b01_011000111000: DATA = 12'b110100100101;
            14'b01_011000111001: DATA = 12'b110100100011;
            14'b01_011000111010: DATA = 12'b110100100001;
            14'b01_011000111011: DATA = 12'b110100011110;
            14'b01_011000111100: DATA = 12'b110100011100;
            14'b01_011000111101: DATA = 12'b110100011001;
            14'b01_011000111110: DATA = 12'b110100010111;
            14'b01_011000111111: DATA = 12'b110100010101;
            14'b01_011001000000: DATA = 12'b110100010010;
            14'b01_011001000001: DATA = 12'b110100010000;
            14'b01_011001000010: DATA = 12'b110100001101;
            14'b01_011001000011: DATA = 12'b110100001011;
            14'b01_011001000100: DATA = 12'b110100001000;
            14'b01_011001000101: DATA = 12'b110100000110;
            14'b01_011001000110: DATA = 12'b110100000011;
            14'b01_011001000111: DATA = 12'b110100000001;
            14'b01_011001001000: DATA = 12'b110011111111;
            14'b01_011001001001: DATA = 12'b110011111100;
            14'b01_011001001010: DATA = 12'b110011111010;
            14'b01_011001001011: DATA = 12'b110011110111;
            14'b01_011001001100: DATA = 12'b110011110101;
            14'b01_011001001101: DATA = 12'b110011110010;
            14'b01_011001001110: DATA = 12'b110011110000;
            14'b01_011001001111: DATA = 12'b110011101101;
            14'b01_011001010000: DATA = 12'b110011101011;
            14'b01_011001010001: DATA = 12'b110011101000;
            14'b01_011001010010: DATA = 12'b110011100110;
            14'b01_011001010011: DATA = 12'b110011100011;
            14'b01_011001010100: DATA = 12'b110011100001;
            14'b01_011001010101: DATA = 12'b110011011110;
            14'b01_011001010110: DATA = 12'b110011011100;
            14'b01_011001010111: DATA = 12'b110011011001;
            14'b01_011001011000: DATA = 12'b110011010111;
            14'b01_011001011001: DATA = 12'b110011010100;
            14'b01_011001011010: DATA = 12'b110011010010;
            14'b01_011001011011: DATA = 12'b110011001111;
            14'b01_011001011100: DATA = 12'b110011001101;
            14'b01_011001011101: DATA = 12'b110011001010;
            14'b01_011001011110: DATA = 12'b110011001000;
            14'b01_011001011111: DATA = 12'b110011000101;
            14'b01_011001100000: DATA = 12'b110011000011;
            14'b01_011001100001: DATA = 12'b110011000000;
            14'b01_011001100010: DATA = 12'b110010111110;
            14'b01_011001100011: DATA = 12'b110010111011;
            14'b01_011001100100: DATA = 12'b110010111001;
            14'b01_011001100101: DATA = 12'b110010110110;
            14'b01_011001100110: DATA = 12'b110010110100;
            14'b01_011001100111: DATA = 12'b110010110001;
            14'b01_011001101000: DATA = 12'b110010101111;
            14'b01_011001101001: DATA = 12'b110010101100;
            14'b01_011001101010: DATA = 12'b110010101010;
            14'b01_011001101011: DATA = 12'b110010100111;
            14'b01_011001101100: DATA = 12'b110010100100;
            14'b01_011001101101: DATA = 12'b110010100010;
            14'b01_011001101110: DATA = 12'b110010011111;
            14'b01_011001101111: DATA = 12'b110010011101;
            14'b01_011001110000: DATA = 12'b110010011010;
            14'b01_011001110001: DATA = 12'b110010011000;
            14'b01_011001110010: DATA = 12'b110010010101;
            14'b01_011001110011: DATA = 12'b110010010010;
            14'b01_011001110100: DATA = 12'b110010010000;
            14'b01_011001110101: DATA = 12'b110010001101;
            14'b01_011001110110: DATA = 12'b110010001011;
            14'b01_011001110111: DATA = 12'b110010001000;
            14'b01_011001111000: DATA = 12'b110010000110;
            14'b01_011001111001: DATA = 12'b110010000011;
            14'b01_011001111010: DATA = 12'b110010000000;
            14'b01_011001111011: DATA = 12'b110001111110;
            14'b01_011001111100: DATA = 12'b110001111011;
            14'b01_011001111101: DATA = 12'b110001111001;
            14'b01_011001111110: DATA = 12'b110001110110;
            14'b01_011001111111: DATA = 12'b110001110011;
            14'b01_011010000000: DATA = 12'b110001110001;
            14'b01_011010000001: DATA = 12'b110001101110;
            14'b01_011010000010: DATA = 12'b110001101100;
            14'b01_011010000011: DATA = 12'b110001101001;
            14'b01_011010000100: DATA = 12'b110001100110;
            14'b01_011010000101: DATA = 12'b110001100100;
            14'b01_011010000110: DATA = 12'b110001100001;
            14'b01_011010000111: DATA = 12'b110001011110;
            14'b01_011010001000: DATA = 12'b110001011100;
            14'b01_011010001001: DATA = 12'b110001011001;
            14'b01_011010001010: DATA = 12'b110001010111;
            14'b01_011010001011: DATA = 12'b110001010100;
            14'b01_011010001100: DATA = 12'b110001010001;
            14'b01_011010001101: DATA = 12'b110001001111;
            14'b01_011010001110: DATA = 12'b110001001100;
            14'b01_011010001111: DATA = 12'b110001001001;
            14'b01_011010010000: DATA = 12'b110001000111;
            14'b01_011010010001: DATA = 12'b110001000100;
            14'b01_011010010010: DATA = 12'b110001000001;
            14'b01_011010010011: DATA = 12'b110000111111;
            14'b01_011010010100: DATA = 12'b110000111100;
            14'b01_011010010101: DATA = 12'b110000111001;
            14'b01_011010010110: DATA = 12'b110000110111;
            14'b01_011010010111: DATA = 12'b110000110100;
            14'b01_011010011000: DATA = 12'b110000110001;
            14'b01_011010011001: DATA = 12'b110000101111;
            14'b01_011010011010: DATA = 12'b110000101100;
            14'b01_011010011011: DATA = 12'b110000101001;
            14'b01_011010011100: DATA = 12'b110000100111;
            14'b01_011010011101: DATA = 12'b110000100100;
            14'b01_011010011110: DATA = 12'b110000100001;
            14'b01_011010011111: DATA = 12'b110000011111;
            14'b01_011010100000: DATA = 12'b110000011100;
            14'b01_011010100001: DATA = 12'b110000011001;
            14'b01_011010100010: DATA = 12'b110000010110;
            14'b01_011010100011: DATA = 12'b110000010100;
            14'b01_011010100100: DATA = 12'b110000010001;
            14'b01_011010100101: DATA = 12'b110000001110;
            14'b01_011010100110: DATA = 12'b110000001100;
            14'b01_011010100111: DATA = 12'b110000001001;
            14'b01_011010101000: DATA = 12'b110000000110;
            14'b01_011010101001: DATA = 12'b110000000100;
            14'b01_011010101010: DATA = 12'b110000000001;
            14'b01_011010101011: DATA = 12'b101111111110;
            14'b01_011010101100: DATA = 12'b101111111011;
            14'b01_011010101101: DATA = 12'b101111111001;
            14'b01_011010101110: DATA = 12'b101111110110;
            14'b01_011010101111: DATA = 12'b101111110011;
            14'b01_011010110000: DATA = 12'b101111110000;
            14'b01_011010110001: DATA = 12'b101111101110;
            14'b01_011010110010: DATA = 12'b101111101011;
            14'b01_011010110011: DATA = 12'b101111101000;
            14'b01_011010110100: DATA = 12'b101111100110;
            14'b01_011010110101: DATA = 12'b101111100011;
            14'b01_011010110110: DATA = 12'b101111100000;
            14'b01_011010110111: DATA = 12'b101111011101;
            14'b01_011010111000: DATA = 12'b101111011011;
            14'b01_011010111001: DATA = 12'b101111011000;
            14'b01_011010111010: DATA = 12'b101111010101;
            14'b01_011010111011: DATA = 12'b101111010010;
            14'b01_011010111100: DATA = 12'b101111010000;
            14'b01_011010111101: DATA = 12'b101111001101;
            14'b01_011010111110: DATA = 12'b101111001010;
            14'b01_011010111111: DATA = 12'b101111000111;
            14'b01_011011000000: DATA = 12'b101111000100;
            14'b01_011011000001: DATA = 12'b101111000010;
            14'b01_011011000010: DATA = 12'b101110111111;
            14'b01_011011000011: DATA = 12'b101110111100;
            14'b01_011011000100: DATA = 12'b101110111001;
            14'b01_011011000101: DATA = 12'b101110110111;
            14'b01_011011000110: DATA = 12'b101110110100;
            14'b01_011011000111: DATA = 12'b101110110001;
            14'b01_011011001000: DATA = 12'b101110101110;
            14'b01_011011001001: DATA = 12'b101110101011;
            14'b01_011011001010: DATA = 12'b101110101001;
            14'b01_011011001011: DATA = 12'b101110100110;
            14'b01_011011001100: DATA = 12'b101110100011;
            14'b01_011011001101: DATA = 12'b101110100000;
            14'b01_011011001110: DATA = 12'b101110011101;
            14'b01_011011001111: DATA = 12'b101110011011;
            14'b01_011011010000: DATA = 12'b101110011000;
            14'b01_011011010001: DATA = 12'b101110010101;
            14'b01_011011010010: DATA = 12'b101110010010;
            14'b01_011011010011: DATA = 12'b101110001111;
            14'b01_011011010100: DATA = 12'b101110001101;
            14'b01_011011010101: DATA = 12'b101110001010;
            14'b01_011011010110: DATA = 12'b101110000111;
            14'b01_011011010111: DATA = 12'b101110000100;
            14'b01_011011011000: DATA = 12'b101110000001;
            14'b01_011011011001: DATA = 12'b101101111111;
            14'b01_011011011010: DATA = 12'b101101111100;
            14'b01_011011011011: DATA = 12'b101101111001;
            14'b01_011011011100: DATA = 12'b101101110110;
            14'b01_011011011101: DATA = 12'b101101110011;
            14'b01_011011011110: DATA = 12'b101101110000;
            14'b01_011011011111: DATA = 12'b101101101110;
            14'b01_011011100000: DATA = 12'b101101101011;
            14'b01_011011100001: DATA = 12'b101101101000;
            14'b01_011011100010: DATA = 12'b101101100101;
            14'b01_011011100011: DATA = 12'b101101100010;
            14'b01_011011100100: DATA = 12'b101101011111;
            14'b01_011011100101: DATA = 12'b101101011100;
            14'b01_011011100110: DATA = 12'b101101011010;
            14'b01_011011100111: DATA = 12'b101101010111;
            14'b01_011011101000: DATA = 12'b101101010100;
            14'b01_011011101001: DATA = 12'b101101010001;
            14'b01_011011101010: DATA = 12'b101101001110;
            14'b01_011011101011: DATA = 12'b101101001011;
            14'b01_011011101100: DATA = 12'b101101001000;
            14'b01_011011101101: DATA = 12'b101101000110;
            14'b01_011011101110: DATA = 12'b101101000011;
            14'b01_011011101111: DATA = 12'b101101000000;
            14'b01_011011110000: DATA = 12'b101100111101;
            14'b01_011011110001: DATA = 12'b101100111010;
            14'b01_011011110010: DATA = 12'b101100110111;
            14'b01_011011110011: DATA = 12'b101100110100;
            14'b01_011011110100: DATA = 12'b101100110010;
            14'b01_011011110101: DATA = 12'b101100101111;
            14'b01_011011110110: DATA = 12'b101100101100;
            14'b01_011011110111: DATA = 12'b101100101001;
            14'b01_011011111000: DATA = 12'b101100100110;
            14'b01_011011111001: DATA = 12'b101100100011;
            14'b01_011011111010: DATA = 12'b101100100000;
            14'b01_011011111011: DATA = 12'b101100011101;
            14'b01_011011111100: DATA = 12'b101100011010;
            14'b01_011011111101: DATA = 12'b101100011000;
            14'b01_011011111110: DATA = 12'b101100010101;
            14'b01_011011111111: DATA = 12'b101100010010;
            14'b01_011100000000: DATA = 12'b101100001111;
            14'b01_011100000001: DATA = 12'b101100001100;
            14'b01_011100000010: DATA = 12'b101100001001;
            14'b01_011100000011: DATA = 12'b101100000110;
            14'b01_011100000100: DATA = 12'b101100000011;
            14'b01_011100000101: DATA = 12'b101100000000;
            14'b01_011100000110: DATA = 12'b101011111101;
            14'b01_011100000111: DATA = 12'b101011111011;
            14'b01_011100001000: DATA = 12'b101011111000;
            14'b01_011100001001: DATA = 12'b101011110101;
            14'b01_011100001010: DATA = 12'b101011110010;
            14'b01_011100001011: DATA = 12'b101011101111;
            14'b01_011100001100: DATA = 12'b101011101100;
            14'b01_011100001101: DATA = 12'b101011101001;
            14'b01_011100001110: DATA = 12'b101011100110;
            14'b01_011100001111: DATA = 12'b101011100011;
            14'b01_011100010000: DATA = 12'b101011100000;
            14'b01_011100010001: DATA = 12'b101011011101;
            14'b01_011100010010: DATA = 12'b101011011010;
            14'b01_011100010011: DATA = 12'b101011010111;
            14'b01_011100010100: DATA = 12'b101011010100;
            14'b01_011100010101: DATA = 12'b101011010010;
            14'b01_011100010110: DATA = 12'b101011001111;
            14'b01_011100010111: DATA = 12'b101011001100;
            14'b01_011100011000: DATA = 12'b101011001001;
            14'b01_011100011001: DATA = 12'b101011000110;
            14'b01_011100011010: DATA = 12'b101011000011;
            14'b01_011100011011: DATA = 12'b101011000000;
            14'b01_011100011100: DATA = 12'b101010111101;
            14'b01_011100011101: DATA = 12'b101010111010;
            14'b01_011100011110: DATA = 12'b101010110111;
            14'b01_011100011111: DATA = 12'b101010110100;
            14'b01_011100100000: DATA = 12'b101010110001;
            14'b01_011100100001: DATA = 12'b101010101110;
            14'b01_011100100010: DATA = 12'b101010101011;
            14'b01_011100100011: DATA = 12'b101010101000;
            14'b01_011100100100: DATA = 12'b101010100101;
            14'b01_011100100101: DATA = 12'b101010100010;
            14'b01_011100100110: DATA = 12'b101010011111;
            14'b01_011100100111: DATA = 12'b101010011100;
            14'b01_011100101000: DATA = 12'b101010011001;
            14'b01_011100101001: DATA = 12'b101010010110;
            14'b01_011100101010: DATA = 12'b101010010011;
            14'b01_011100101011: DATA = 12'b101010010000;
            14'b01_011100101100: DATA = 12'b101010001110;
            14'b01_011100101101: DATA = 12'b101010001011;
            14'b01_011100101110: DATA = 12'b101010001000;
            14'b01_011100101111: DATA = 12'b101010000101;
            14'b01_011100110000: DATA = 12'b101010000010;
            14'b01_011100110001: DATA = 12'b101001111111;
            14'b01_011100110010: DATA = 12'b101001111100;
            14'b01_011100110011: DATA = 12'b101001111001;
            14'b01_011100110100: DATA = 12'b101001110110;
            14'b01_011100110101: DATA = 12'b101001110011;
            14'b01_011100110110: DATA = 12'b101001110000;
            14'b01_011100110111: DATA = 12'b101001101101;
            14'b01_011100111000: DATA = 12'b101001101010;
            14'b01_011100111001: DATA = 12'b101001100111;
            14'b01_011100111010: DATA = 12'b101001100100;
            14'b01_011100111011: DATA = 12'b101001100001;
            14'b01_011100111100: DATA = 12'b101001011110;
            14'b01_011100111101: DATA = 12'b101001011011;
            14'b01_011100111110: DATA = 12'b101001011000;
            14'b01_011100111111: DATA = 12'b101001010101;
            14'b01_011101000000: DATA = 12'b101001010010;
            14'b01_011101000001: DATA = 12'b101001001111;
            14'b01_011101000010: DATA = 12'b101001001100;
            14'b01_011101000011: DATA = 12'b101001001001;
            14'b01_011101000100: DATA = 12'b101001000110;
            14'b01_011101000101: DATA = 12'b101001000011;
            14'b01_011101000110: DATA = 12'b101001000000;
            14'b01_011101000111: DATA = 12'b101000111101;
            14'b01_011101001000: DATA = 12'b101000111010;
            14'b01_011101001001: DATA = 12'b101000110111;
            14'b01_011101001010: DATA = 12'b101000110100;
            14'b01_011101001011: DATA = 12'b101000110001;
            14'b01_011101001100: DATA = 12'b101000101110;
            14'b01_011101001101: DATA = 12'b101000101011;
            14'b01_011101001110: DATA = 12'b101000101000;
            14'b01_011101001111: DATA = 12'b101000100100;
            14'b01_011101010000: DATA = 12'b101000100001;
            14'b01_011101010001: DATA = 12'b101000011110;
            14'b01_011101010010: DATA = 12'b101000011011;
            14'b01_011101010011: DATA = 12'b101000011000;
            14'b01_011101010100: DATA = 12'b101000010101;
            14'b01_011101010101: DATA = 12'b101000010010;
            14'b01_011101010110: DATA = 12'b101000001111;
            14'b01_011101010111: DATA = 12'b101000001100;
            14'b01_011101011000: DATA = 12'b101000001001;
            14'b01_011101011001: DATA = 12'b101000000110;
            14'b01_011101011010: DATA = 12'b101000000011;
            14'b01_011101011011: DATA = 12'b101000000000;
            14'b01_011101011100: DATA = 12'b100111111101;
            14'b01_011101011101: DATA = 12'b100111111010;
            14'b01_011101011110: DATA = 12'b100111110111;
            14'b01_011101011111: DATA = 12'b100111110100;
            14'b01_011101100000: DATA = 12'b100111110001;
            14'b01_011101100001: DATA = 12'b100111101110;
            14'b01_011101100010: DATA = 12'b100111101011;
            14'b01_011101100011: DATA = 12'b100111101000;
            14'b01_011101100100: DATA = 12'b100111100101;
            14'b01_011101100101: DATA = 12'b100111100010;
            14'b01_011101100110: DATA = 12'b100111011111;
            14'b01_011101100111: DATA = 12'b100111011100;
            14'b01_011101101000: DATA = 12'b100111011000;
            14'b01_011101101001: DATA = 12'b100111010101;
            14'b01_011101101010: DATA = 12'b100111010010;
            14'b01_011101101011: DATA = 12'b100111001111;
            14'b01_011101101100: DATA = 12'b100111001100;
            14'b01_011101101101: DATA = 12'b100111001001;
            14'b01_011101101110: DATA = 12'b100111000110;
            14'b01_011101101111: DATA = 12'b100111000011;
            14'b01_011101110000: DATA = 12'b100111000000;
            14'b01_011101110001: DATA = 12'b100110111101;
            14'b01_011101110010: DATA = 12'b100110111010;
            14'b01_011101110011: DATA = 12'b100110110111;
            14'b01_011101110100: DATA = 12'b100110110100;
            14'b01_011101110101: DATA = 12'b100110110001;
            14'b01_011101110110: DATA = 12'b100110101110;
            14'b01_011101110111: DATA = 12'b100110101011;
            14'b01_011101111000: DATA = 12'b100110100111;
            14'b01_011101111001: DATA = 12'b100110100100;
            14'b01_011101111010: DATA = 12'b100110100001;
            14'b01_011101111011: DATA = 12'b100110011110;
            14'b01_011101111100: DATA = 12'b100110011011;
            14'b01_011101111101: DATA = 12'b100110011000;
            14'b01_011101111110: DATA = 12'b100110010101;
            14'b01_011101111111: DATA = 12'b100110010010;
            14'b01_011110000000: DATA = 12'b100110001111;
            14'b01_011110000001: DATA = 12'b100110001100;
            14'b01_011110000010: DATA = 12'b100110001001;
            14'b01_011110000011: DATA = 12'b100110000110;
            14'b01_011110000100: DATA = 12'b100110000011;
            14'b01_011110000101: DATA = 12'b100101111111;
            14'b01_011110000110: DATA = 12'b100101111100;
            14'b01_011110000111: DATA = 12'b100101111001;
            14'b01_011110001000: DATA = 12'b100101110110;
            14'b01_011110001001: DATA = 12'b100101110011;
            14'b01_011110001010: DATA = 12'b100101110000;
            14'b01_011110001011: DATA = 12'b100101101101;
            14'b01_011110001100: DATA = 12'b100101101010;
            14'b01_011110001101: DATA = 12'b100101100111;
            14'b01_011110001110: DATA = 12'b100101100100;
            14'b01_011110001111: DATA = 12'b100101100001;
            14'b01_011110010000: DATA = 12'b100101011101;
            14'b01_011110010001: DATA = 12'b100101011010;
            14'b01_011110010010: DATA = 12'b100101010111;
            14'b01_011110010011: DATA = 12'b100101010100;
            14'b01_011110010100: DATA = 12'b100101010001;
            14'b01_011110010101: DATA = 12'b100101001110;
            14'b01_011110010110: DATA = 12'b100101001011;
            14'b01_011110010111: DATA = 12'b100101001000;
            14'b01_011110011000: DATA = 12'b100101000101;
            14'b01_011110011001: DATA = 12'b100101000010;
            14'b01_011110011010: DATA = 12'b100100111110;
            14'b01_011110011011: DATA = 12'b100100111011;
            14'b01_011110011100: DATA = 12'b100100111000;
            14'b01_011110011101: DATA = 12'b100100110101;
            14'b01_011110011110: DATA = 12'b100100110010;
            14'b01_011110011111: DATA = 12'b100100101111;
            14'b01_011110100000: DATA = 12'b100100101100;
            14'b01_011110100001: DATA = 12'b100100101001;
            14'b01_011110100010: DATA = 12'b100100100110;
            14'b01_011110100011: DATA = 12'b100100100011;
            14'b01_011110100100: DATA = 12'b100100011111;
            14'b01_011110100101: DATA = 12'b100100011100;
            14'b01_011110100110: DATA = 12'b100100011001;
            14'b01_011110100111: DATA = 12'b100100010110;
            14'b01_011110101000: DATA = 12'b100100010011;
            14'b01_011110101001: DATA = 12'b100100010000;
            14'b01_011110101010: DATA = 12'b100100001101;
            14'b01_011110101011: DATA = 12'b100100001010;
            14'b01_011110101100: DATA = 12'b100100000111;
            14'b01_011110101101: DATA = 12'b100100000011;
            14'b01_011110101110: DATA = 12'b100100000000;
            14'b01_011110101111: DATA = 12'b100011111101;
            14'b01_011110110000: DATA = 12'b100011111010;
            14'b01_011110110001: DATA = 12'b100011110111;
            14'b01_011110110010: DATA = 12'b100011110100;
            14'b01_011110110011: DATA = 12'b100011110001;
            14'b01_011110110100: DATA = 12'b100011101110;
            14'b01_011110110101: DATA = 12'b100011101010;
            14'b01_011110110110: DATA = 12'b100011100111;
            14'b01_011110110111: DATA = 12'b100011100100;
            14'b01_011110111000: DATA = 12'b100011100001;
            14'b01_011110111001: DATA = 12'b100011011110;
            14'b01_011110111010: DATA = 12'b100011011011;
            14'b01_011110111011: DATA = 12'b100011011000;
            14'b01_011110111100: DATA = 12'b100011010101;
            14'b01_011110111101: DATA = 12'b100011010010;
            14'b01_011110111110: DATA = 12'b100011001110;
            14'b01_011110111111: DATA = 12'b100011001011;
            14'b01_011111000000: DATA = 12'b100011001000;
            14'b01_011111000001: DATA = 12'b100011000101;
            14'b01_011111000010: DATA = 12'b100011000010;
            14'b01_011111000011: DATA = 12'b100010111111;
            14'b01_011111000100: DATA = 12'b100010111100;
            14'b01_011111000101: DATA = 12'b100010111001;
            14'b01_011111000110: DATA = 12'b100010110101;
            14'b01_011111000111: DATA = 12'b100010110010;
            14'b01_011111001000: DATA = 12'b100010101111;
            14'b01_011111001001: DATA = 12'b100010101100;
            14'b01_011111001010: DATA = 12'b100010101001;
            14'b01_011111001011: DATA = 12'b100010100110;
            14'b01_011111001100: DATA = 12'b100010100011;
            14'b01_011111001101: DATA = 12'b100010011111;
            14'b01_011111001110: DATA = 12'b100010011100;
            14'b01_011111001111: DATA = 12'b100010011001;
            14'b01_011111010000: DATA = 12'b100010010110;
            14'b01_011111010001: DATA = 12'b100010010011;
            14'b01_011111010010: DATA = 12'b100010010000;
            14'b01_011111010011: DATA = 12'b100010001101;
            14'b01_011111010100: DATA = 12'b100010001010;
            14'b01_011111010101: DATA = 12'b100010000110;
            14'b01_011111010110: DATA = 12'b100010000011;
            14'b01_011111010111: DATA = 12'b100010000000;
            14'b01_011111011000: DATA = 12'b100001111101;
            14'b01_011111011001: DATA = 12'b100001111010;
            14'b01_011111011010: DATA = 12'b100001110111;
            14'b01_011111011011: DATA = 12'b100001110100;
            14'b01_011111011100: DATA = 12'b100001110000;
            14'b01_011111011101: DATA = 12'b100001101101;
            14'b01_011111011110: DATA = 12'b100001101010;
            14'b01_011111011111: DATA = 12'b100001100111;
            14'b01_011111100000: DATA = 12'b100001100100;
            14'b01_011111100001: DATA = 12'b100001100001;
            14'b01_011111100010: DATA = 12'b100001011110;
            14'b01_011111100011: DATA = 12'b100001011011;
            14'b01_011111100100: DATA = 12'b100001010111;
            14'b01_011111100101: DATA = 12'b100001010100;
            14'b01_011111100110: DATA = 12'b100001010001;
            14'b01_011111100111: DATA = 12'b100001001110;
            14'b01_011111101000: DATA = 12'b100001001011;
            14'b01_011111101001: DATA = 12'b100001001000;
            14'b01_011111101010: DATA = 12'b100001000101;
            14'b01_011111101011: DATA = 12'b100001000001;
            14'b01_011111101100: DATA = 12'b100000111110;
            14'b01_011111101101: DATA = 12'b100000111011;
            14'b01_011111101110: DATA = 12'b100000111000;
            14'b01_011111101111: DATA = 12'b100000110101;
            14'b01_011111110000: DATA = 12'b100000110010;
            14'b01_011111110001: DATA = 12'b100000101111;
            14'b01_011111110010: DATA = 12'b100000101011;
            14'b01_011111110011: DATA = 12'b100000101000;
            14'b01_011111110100: DATA = 12'b100000100101;
            14'b01_011111110101: DATA = 12'b100000100010;
            14'b01_011111110110: DATA = 12'b100000011111;
            14'b01_011111110111: DATA = 12'b100000011100;
            14'b01_011111111000: DATA = 12'b100000011001;
            14'b01_011111111001: DATA = 12'b100000010101;
            14'b01_011111111010: DATA = 12'b100000010010;
            14'b01_011111111011: DATA = 12'b100000001111;
            14'b01_011111111100: DATA = 12'b100000001100;
            14'b01_011111111101: DATA = 12'b100000001001;
            14'b01_011111111110: DATA = 12'b100000000110;
            14'b01_011111111111: DATA = 12'b100000000011;
            14'b01_100000000000: DATA = 12'b100000000000;
            14'b01_100000000001: DATA = 12'b100000000000;
            14'b01_100000000010: DATA = 12'b100000000000;
            14'b01_100000000011: DATA = 12'b100000000000;
            14'b01_100000000100: DATA = 12'b100000000000;
            14'b01_100000000101: DATA = 12'b100000000000;
            14'b01_100000000110: DATA = 12'b100000000000;
            14'b01_100000000111: DATA = 12'b100000000000;
            14'b01_100000001000: DATA = 12'b100000000000;
            14'b01_100000001001: DATA = 12'b100000000000;
            14'b01_100000001010: DATA = 12'b100000000000;
            14'b01_100000001011: DATA = 12'b100000000000;
            14'b01_100000001100: DATA = 12'b100000000000;
            14'b01_100000001101: DATA = 12'b100000000000;
            14'b01_100000001110: DATA = 12'b100000000000;
            14'b01_100000001111: DATA = 12'b100000000000;
            14'b01_100000010000: DATA = 12'b100000000000;
            14'b01_100000010001: DATA = 12'b100000000000;
            14'b01_100000010010: DATA = 12'b100000000000;
            14'b01_100000010011: DATA = 12'b100000000000;
            14'b01_100000010100: DATA = 12'b100000000000;
            14'b01_100000010101: DATA = 12'b100000000000;
            14'b01_100000010110: DATA = 12'b100000000000;
            14'b01_100000010111: DATA = 12'b100000000000;
            14'b01_100000011000: DATA = 12'b100000000000;
            14'b01_100000011001: DATA = 12'b100000000000;
            14'b01_100000011010: DATA = 12'b100000000000;
            14'b01_100000011011: DATA = 12'b100000000000;
            14'b01_100000011100: DATA = 12'b100000000000;
            14'b01_100000011101: DATA = 12'b100000000000;
            14'b01_100000011110: DATA = 12'b100000000000;
            14'b01_100000011111: DATA = 12'b100000000000;
            14'b01_100000100000: DATA = 12'b100000000000;
            14'b01_100000100001: DATA = 12'b100000000000;
            14'b01_100000100010: DATA = 12'b100000000000;
            14'b01_100000100011: DATA = 12'b100000000000;
            14'b01_100000100100: DATA = 12'b100000000000;
            14'b01_100000100101: DATA = 12'b100000000000;
            14'b01_100000100110: DATA = 12'b100000000000;
            14'b01_100000100111: DATA = 12'b100000000000;
            14'b01_100000101000: DATA = 12'b100000000000;
            14'b01_100000101001: DATA = 12'b100000000000;
            14'b01_100000101010: DATA = 12'b100000000000;
            14'b01_100000101011: DATA = 12'b100000000000;
            14'b01_100000101100: DATA = 12'b100000000000;
            14'b01_100000101101: DATA = 12'b100000000000;
            14'b01_100000101110: DATA = 12'b100000000000;
            14'b01_100000101111: DATA = 12'b100000000000;
            14'b01_100000110000: DATA = 12'b100000000000;
            14'b01_100000110001: DATA = 12'b100000000000;
            14'b01_100000110010: DATA = 12'b100000000000;
            14'b01_100000110011: DATA = 12'b100000000000;
            14'b01_100000110100: DATA = 12'b100000000000;
            14'b01_100000110101: DATA = 12'b100000000000;
            14'b01_100000110110: DATA = 12'b100000000000;
            14'b01_100000110111: DATA = 12'b100000000000;
            14'b01_100000111000: DATA = 12'b100000000000;
            14'b01_100000111001: DATA = 12'b100000000000;
            14'b01_100000111010: DATA = 12'b100000000000;
            14'b01_100000111011: DATA = 12'b100000000000;
            14'b01_100000111100: DATA = 12'b100000000000;
            14'b01_100000111101: DATA = 12'b100000000000;
            14'b01_100000111110: DATA = 12'b100000000000;
            14'b01_100000111111: DATA = 12'b100000000000;
            14'b01_100001000000: DATA = 12'b100000000000;
            14'b01_100001000001: DATA = 12'b100000000000;
            14'b01_100001000010: DATA = 12'b100000000000;
            14'b01_100001000011: DATA = 12'b100000000000;
            14'b01_100001000100: DATA = 12'b100000000000;
            14'b01_100001000101: DATA = 12'b100000000000;
            14'b01_100001000110: DATA = 12'b100000000000;
            14'b01_100001000111: DATA = 12'b100000000000;
            14'b01_100001001000: DATA = 12'b100000000000;
            14'b01_100001001001: DATA = 12'b100000000000;
            14'b01_100001001010: DATA = 12'b100000000000;
            14'b01_100001001011: DATA = 12'b100000000000;
            14'b01_100001001100: DATA = 12'b100000000000;
            14'b01_100001001101: DATA = 12'b100000000000;
            14'b01_100001001110: DATA = 12'b100000000000;
            14'b01_100001001111: DATA = 12'b100000000000;
            14'b01_100001010000: DATA = 12'b100000000000;
            14'b01_100001010001: DATA = 12'b100000000000;
            14'b01_100001010010: DATA = 12'b100000000000;
            14'b01_100001010011: DATA = 12'b100000000000;
            14'b01_100001010100: DATA = 12'b100000000000;
            14'b01_100001010101: DATA = 12'b100000000000;
            14'b01_100001010110: DATA = 12'b100000000000;
            14'b01_100001010111: DATA = 12'b100000000000;
            14'b01_100001011000: DATA = 12'b100000000000;
            14'b01_100001011001: DATA = 12'b100000000000;
            14'b01_100001011010: DATA = 12'b100000000000;
            14'b01_100001011011: DATA = 12'b100000000000;
            14'b01_100001011100: DATA = 12'b100000000000;
            14'b01_100001011101: DATA = 12'b100000000000;
            14'b01_100001011110: DATA = 12'b100000000000;
            14'b01_100001011111: DATA = 12'b100000000000;
            14'b01_100001100000: DATA = 12'b100000000000;
            14'b01_100001100001: DATA = 12'b100000000000;
            14'b01_100001100010: DATA = 12'b100000000000;
            14'b01_100001100011: DATA = 12'b100000000000;
            14'b01_100001100100: DATA = 12'b100000000000;
            14'b01_100001100101: DATA = 12'b100000000000;
            14'b01_100001100110: DATA = 12'b100000000000;
            14'b01_100001100111: DATA = 12'b100000000000;
            14'b01_100001101000: DATA = 12'b100000000000;
            14'b01_100001101001: DATA = 12'b100000000000;
            14'b01_100001101010: DATA = 12'b100000000000;
            14'b01_100001101011: DATA = 12'b100000000000;
            14'b01_100001101100: DATA = 12'b100000000000;
            14'b01_100001101101: DATA = 12'b100000000000;
            14'b01_100001101110: DATA = 12'b100000000000;
            14'b01_100001101111: DATA = 12'b100000000000;
            14'b01_100001110000: DATA = 12'b100000000000;
            14'b01_100001110001: DATA = 12'b100000000000;
            14'b01_100001110010: DATA = 12'b100000000000;
            14'b01_100001110011: DATA = 12'b100000000000;
            14'b01_100001110100: DATA = 12'b100000000000;
            14'b01_100001110101: DATA = 12'b100000000000;
            14'b01_100001110110: DATA = 12'b100000000000;
            14'b01_100001110111: DATA = 12'b100000000000;
            14'b01_100001111000: DATA = 12'b100000000000;
            14'b01_100001111001: DATA = 12'b100000000000;
            14'b01_100001111010: DATA = 12'b100000000000;
            14'b01_100001111011: DATA = 12'b100000000000;
            14'b01_100001111100: DATA = 12'b100000000000;
            14'b01_100001111101: DATA = 12'b100000000000;
            14'b01_100001111110: DATA = 12'b100000000000;
            14'b01_100001111111: DATA = 12'b100000000000;
            14'b01_100010000000: DATA = 12'b100000000000;
            14'b01_100010000001: DATA = 12'b100000000000;
            14'b01_100010000010: DATA = 12'b100000000000;
            14'b01_100010000011: DATA = 12'b100000000000;
            14'b01_100010000100: DATA = 12'b100000000000;
            14'b01_100010000101: DATA = 12'b100000000000;
            14'b01_100010000110: DATA = 12'b100000000000;
            14'b01_100010000111: DATA = 12'b100000000000;
            14'b01_100010001000: DATA = 12'b100000000000;
            14'b01_100010001001: DATA = 12'b100000000000;
            14'b01_100010001010: DATA = 12'b100000000000;
            14'b01_100010001011: DATA = 12'b100000000000;
            14'b01_100010001100: DATA = 12'b100000000000;
            14'b01_100010001101: DATA = 12'b100000000000;
            14'b01_100010001110: DATA = 12'b100000000000;
            14'b01_100010001111: DATA = 12'b100000000000;
            14'b01_100010010000: DATA = 12'b100000000000;
            14'b01_100010010001: DATA = 12'b100000000000;
            14'b01_100010010010: DATA = 12'b100000000000;
            14'b01_100010010011: DATA = 12'b100000000000;
            14'b01_100010010100: DATA = 12'b100000000000;
            14'b01_100010010101: DATA = 12'b100000000000;
            14'b01_100010010110: DATA = 12'b100000000000;
            14'b01_100010010111: DATA = 12'b100000000000;
            14'b01_100010011000: DATA = 12'b100000000000;
            14'b01_100010011001: DATA = 12'b100000000000;
            14'b01_100010011010: DATA = 12'b100000000000;
            14'b01_100010011011: DATA = 12'b100000000000;
            14'b01_100010011100: DATA = 12'b100000000000;
            14'b01_100010011101: DATA = 12'b100000000000;
            14'b01_100010011110: DATA = 12'b100000000000;
            14'b01_100010011111: DATA = 12'b100000000000;
            14'b01_100010100000: DATA = 12'b100000000000;
            14'b01_100010100001: DATA = 12'b100000000000;
            14'b01_100010100010: DATA = 12'b100000000000;
            14'b01_100010100011: DATA = 12'b100000000000;
            14'b01_100010100100: DATA = 12'b100000000000;
            14'b01_100010100101: DATA = 12'b100000000000;
            14'b01_100010100110: DATA = 12'b100000000000;
            14'b01_100010100111: DATA = 12'b100000000000;
            14'b01_100010101000: DATA = 12'b100000000000;
            14'b01_100010101001: DATA = 12'b100000000000;
            14'b01_100010101010: DATA = 12'b100000000000;
            14'b01_100010101011: DATA = 12'b100000000000;
            14'b01_100010101100: DATA = 12'b100000000000;
            14'b01_100010101101: DATA = 12'b100000000000;
            14'b01_100010101110: DATA = 12'b100000000000;
            14'b01_100010101111: DATA = 12'b100000000000;
            14'b01_100010110000: DATA = 12'b100000000000;
            14'b01_100010110001: DATA = 12'b100000000000;
            14'b01_100010110010: DATA = 12'b100000000000;
            14'b01_100010110011: DATA = 12'b100000000000;
            14'b01_100010110100: DATA = 12'b100000000000;
            14'b01_100010110101: DATA = 12'b100000000000;
            14'b01_100010110110: DATA = 12'b100000000000;
            14'b01_100010110111: DATA = 12'b100000000000;
            14'b01_100010111000: DATA = 12'b100000000000;
            14'b01_100010111001: DATA = 12'b100000000000;
            14'b01_100010111010: DATA = 12'b100000000000;
            14'b01_100010111011: DATA = 12'b100000000000;
            14'b01_100010111100: DATA = 12'b100000000000;
            14'b01_100010111101: DATA = 12'b100000000000;
            14'b01_100010111110: DATA = 12'b100000000000;
            14'b01_100010111111: DATA = 12'b100000000000;
            14'b01_100011000000: DATA = 12'b100000000000;
            14'b01_100011000001: DATA = 12'b100000000000;
            14'b01_100011000010: DATA = 12'b100000000000;
            14'b01_100011000011: DATA = 12'b100000000000;
            14'b01_100011000100: DATA = 12'b100000000000;
            14'b01_100011000101: DATA = 12'b100000000000;
            14'b01_100011000110: DATA = 12'b100000000000;
            14'b01_100011000111: DATA = 12'b100000000000;
            14'b01_100011001000: DATA = 12'b100000000000;
            14'b01_100011001001: DATA = 12'b100000000000;
            14'b01_100011001010: DATA = 12'b100000000000;
            14'b01_100011001011: DATA = 12'b100000000000;
            14'b01_100011001100: DATA = 12'b100000000000;
            14'b01_100011001101: DATA = 12'b100000000000;
            14'b01_100011001110: DATA = 12'b100000000000;
            14'b01_100011001111: DATA = 12'b100000000000;
            14'b01_100011010000: DATA = 12'b100000000000;
            14'b01_100011010001: DATA = 12'b100000000000;
            14'b01_100011010010: DATA = 12'b100000000000;
            14'b01_100011010011: DATA = 12'b100000000000;
            14'b01_100011010100: DATA = 12'b100000000000;
            14'b01_100011010101: DATA = 12'b100000000000;
            14'b01_100011010110: DATA = 12'b100000000000;
            14'b01_100011010111: DATA = 12'b100000000000;
            14'b01_100011011000: DATA = 12'b100000000000;
            14'b01_100011011001: DATA = 12'b100000000000;
            14'b01_100011011010: DATA = 12'b100000000000;
            14'b01_100011011011: DATA = 12'b100000000000;
            14'b01_100011011100: DATA = 12'b100000000000;
            14'b01_100011011101: DATA = 12'b100000000000;
            14'b01_100011011110: DATA = 12'b100000000000;
            14'b01_100011011111: DATA = 12'b100000000000;
            14'b01_100011100000: DATA = 12'b100000000000;
            14'b01_100011100001: DATA = 12'b100000000000;
            14'b01_100011100010: DATA = 12'b100000000000;
            14'b01_100011100011: DATA = 12'b100000000000;
            14'b01_100011100100: DATA = 12'b100000000000;
            14'b01_100011100101: DATA = 12'b100000000000;
            14'b01_100011100110: DATA = 12'b100000000000;
            14'b01_100011100111: DATA = 12'b100000000000;
            14'b01_100011101000: DATA = 12'b100000000000;
            14'b01_100011101001: DATA = 12'b100000000000;
            14'b01_100011101010: DATA = 12'b100000000000;
            14'b01_100011101011: DATA = 12'b100000000000;
            14'b01_100011101100: DATA = 12'b100000000000;
            14'b01_100011101101: DATA = 12'b100000000000;
            14'b01_100011101110: DATA = 12'b100000000000;
            14'b01_100011101111: DATA = 12'b100000000000;
            14'b01_100011110000: DATA = 12'b100000000000;
            14'b01_100011110001: DATA = 12'b100000000000;
            14'b01_100011110010: DATA = 12'b100000000000;
            14'b01_100011110011: DATA = 12'b100000000000;
            14'b01_100011110100: DATA = 12'b100000000000;
            14'b01_100011110101: DATA = 12'b100000000000;
            14'b01_100011110110: DATA = 12'b100000000000;
            14'b01_100011110111: DATA = 12'b100000000000;
            14'b01_100011111000: DATA = 12'b100000000000;
            14'b01_100011111001: DATA = 12'b100000000000;
            14'b01_100011111010: DATA = 12'b100000000000;
            14'b01_100011111011: DATA = 12'b100000000000;
            14'b01_100011111100: DATA = 12'b100000000000;
            14'b01_100011111101: DATA = 12'b100000000000;
            14'b01_100011111110: DATA = 12'b100000000000;
            14'b01_100011111111: DATA = 12'b100000000000;
            14'b01_100100000000: DATA = 12'b100000000000;
            14'b01_100100000001: DATA = 12'b100000000000;
            14'b01_100100000010: DATA = 12'b100000000000;
            14'b01_100100000011: DATA = 12'b100000000000;
            14'b01_100100000100: DATA = 12'b100000000000;
            14'b01_100100000101: DATA = 12'b100000000000;
            14'b01_100100000110: DATA = 12'b100000000000;
            14'b01_100100000111: DATA = 12'b100000000000;
            14'b01_100100001000: DATA = 12'b100000000000;
            14'b01_100100001001: DATA = 12'b100000000000;
            14'b01_100100001010: DATA = 12'b100000000000;
            14'b01_100100001011: DATA = 12'b100000000000;
            14'b01_100100001100: DATA = 12'b100000000000;
            14'b01_100100001101: DATA = 12'b100000000000;
            14'b01_100100001110: DATA = 12'b100000000000;
            14'b01_100100001111: DATA = 12'b100000000000;
            14'b01_100100010000: DATA = 12'b100000000000;
            14'b01_100100010001: DATA = 12'b100000000000;
            14'b01_100100010010: DATA = 12'b100000000000;
            14'b01_100100010011: DATA = 12'b100000000000;
            14'b01_100100010100: DATA = 12'b100000000000;
            14'b01_100100010101: DATA = 12'b100000000000;
            14'b01_100100010110: DATA = 12'b100000000000;
            14'b01_100100010111: DATA = 12'b100000000000;
            14'b01_100100011000: DATA = 12'b100000000000;
            14'b01_100100011001: DATA = 12'b100000000000;
            14'b01_100100011010: DATA = 12'b100000000000;
            14'b01_100100011011: DATA = 12'b100000000000;
            14'b01_100100011100: DATA = 12'b100000000000;
            14'b01_100100011101: DATA = 12'b100000000000;
            14'b01_100100011110: DATA = 12'b100000000000;
            14'b01_100100011111: DATA = 12'b100000000000;
            14'b01_100100100000: DATA = 12'b100000000000;
            14'b01_100100100001: DATA = 12'b100000000000;
            14'b01_100100100010: DATA = 12'b100000000000;
            14'b01_100100100011: DATA = 12'b100000000000;
            14'b01_100100100100: DATA = 12'b100000000000;
            14'b01_100100100101: DATA = 12'b100000000000;
            14'b01_100100100110: DATA = 12'b100000000000;
            14'b01_100100100111: DATA = 12'b100000000000;
            14'b01_100100101000: DATA = 12'b100000000000;
            14'b01_100100101001: DATA = 12'b100000000000;
            14'b01_100100101010: DATA = 12'b100000000000;
            14'b01_100100101011: DATA = 12'b100000000000;
            14'b01_100100101100: DATA = 12'b100000000000;
            14'b01_100100101101: DATA = 12'b100000000000;
            14'b01_100100101110: DATA = 12'b100000000000;
            14'b01_100100101111: DATA = 12'b100000000000;
            14'b01_100100110000: DATA = 12'b100000000000;
            14'b01_100100110001: DATA = 12'b100000000000;
            14'b01_100100110010: DATA = 12'b100000000000;
            14'b01_100100110011: DATA = 12'b100000000000;
            14'b01_100100110100: DATA = 12'b100000000000;
            14'b01_100100110101: DATA = 12'b100000000000;
            14'b01_100100110110: DATA = 12'b100000000000;
            14'b01_100100110111: DATA = 12'b100000000000;
            14'b01_100100111000: DATA = 12'b100000000000;
            14'b01_100100111001: DATA = 12'b100000000000;
            14'b01_100100111010: DATA = 12'b100000000000;
            14'b01_100100111011: DATA = 12'b100000000000;
            14'b01_100100111100: DATA = 12'b100000000000;
            14'b01_100100111101: DATA = 12'b100000000000;
            14'b01_100100111110: DATA = 12'b100000000000;
            14'b01_100100111111: DATA = 12'b100000000000;
            14'b01_100101000000: DATA = 12'b100000000000;
            14'b01_100101000001: DATA = 12'b100000000000;
            14'b01_100101000010: DATA = 12'b100000000000;
            14'b01_100101000011: DATA = 12'b100000000000;
            14'b01_100101000100: DATA = 12'b100000000000;
            14'b01_100101000101: DATA = 12'b100000000000;
            14'b01_100101000110: DATA = 12'b100000000000;
            14'b01_100101000111: DATA = 12'b100000000000;
            14'b01_100101001000: DATA = 12'b100000000000;
            14'b01_100101001001: DATA = 12'b100000000000;
            14'b01_100101001010: DATA = 12'b100000000000;
            14'b01_100101001011: DATA = 12'b100000000000;
            14'b01_100101001100: DATA = 12'b100000000000;
            14'b01_100101001101: DATA = 12'b100000000000;
            14'b01_100101001110: DATA = 12'b100000000000;
            14'b01_100101001111: DATA = 12'b100000000000;
            14'b01_100101010000: DATA = 12'b100000000000;
            14'b01_100101010001: DATA = 12'b100000000000;
            14'b01_100101010010: DATA = 12'b100000000000;
            14'b01_100101010011: DATA = 12'b100000000000;
            14'b01_100101010100: DATA = 12'b100000000000;
            14'b01_100101010101: DATA = 12'b100000000000;
            14'b01_100101010110: DATA = 12'b100000000000;
            14'b01_100101010111: DATA = 12'b100000000000;
            14'b01_100101011000: DATA = 12'b100000000000;
            14'b01_100101011001: DATA = 12'b100000000000;
            14'b01_100101011010: DATA = 12'b100000000000;
            14'b01_100101011011: DATA = 12'b100000000000;
            14'b01_100101011100: DATA = 12'b100000000000;
            14'b01_100101011101: DATA = 12'b100000000000;
            14'b01_100101011110: DATA = 12'b100000000000;
            14'b01_100101011111: DATA = 12'b100000000000;
            14'b01_100101100000: DATA = 12'b100000000000;
            14'b01_100101100001: DATA = 12'b100000000000;
            14'b01_100101100010: DATA = 12'b100000000000;
            14'b01_100101100011: DATA = 12'b100000000000;
            14'b01_100101100100: DATA = 12'b100000000000;
            14'b01_100101100101: DATA = 12'b100000000000;
            14'b01_100101100110: DATA = 12'b100000000000;
            14'b01_100101100111: DATA = 12'b100000000000;
            14'b01_100101101000: DATA = 12'b100000000000;
            14'b01_100101101001: DATA = 12'b100000000000;
            14'b01_100101101010: DATA = 12'b100000000000;
            14'b01_100101101011: DATA = 12'b100000000000;
            14'b01_100101101100: DATA = 12'b100000000000;
            14'b01_100101101101: DATA = 12'b100000000000;
            14'b01_100101101110: DATA = 12'b100000000000;
            14'b01_100101101111: DATA = 12'b100000000000;
            14'b01_100101110000: DATA = 12'b100000000000;
            14'b01_100101110001: DATA = 12'b100000000000;
            14'b01_100101110010: DATA = 12'b100000000000;
            14'b01_100101110011: DATA = 12'b100000000000;
            14'b01_100101110100: DATA = 12'b100000000000;
            14'b01_100101110101: DATA = 12'b100000000000;
            14'b01_100101110110: DATA = 12'b100000000000;
            14'b01_100101110111: DATA = 12'b100000000000;
            14'b01_100101111000: DATA = 12'b100000000000;
            14'b01_100101111001: DATA = 12'b100000000000;
            14'b01_100101111010: DATA = 12'b100000000000;
            14'b01_100101111011: DATA = 12'b100000000000;
            14'b01_100101111100: DATA = 12'b100000000000;
            14'b01_100101111101: DATA = 12'b100000000000;
            14'b01_100101111110: DATA = 12'b100000000000;
            14'b01_100101111111: DATA = 12'b100000000000;
            14'b01_100110000000: DATA = 12'b100000000000;
            14'b01_100110000001: DATA = 12'b100000000000;
            14'b01_100110000010: DATA = 12'b100000000000;
            14'b01_100110000011: DATA = 12'b100000000000;
            14'b01_100110000100: DATA = 12'b100000000000;
            14'b01_100110000101: DATA = 12'b100000000000;
            14'b01_100110000110: DATA = 12'b100000000000;
            14'b01_100110000111: DATA = 12'b100000000000;
            14'b01_100110001000: DATA = 12'b100000000000;
            14'b01_100110001001: DATA = 12'b100000000000;
            14'b01_100110001010: DATA = 12'b100000000000;
            14'b01_100110001011: DATA = 12'b100000000000;
            14'b01_100110001100: DATA = 12'b100000000000;
            14'b01_100110001101: DATA = 12'b100000000000;
            14'b01_100110001110: DATA = 12'b100000000000;
            14'b01_100110001111: DATA = 12'b100000000000;
            14'b01_100110010000: DATA = 12'b100000000000;
            14'b01_100110010001: DATA = 12'b100000000000;
            14'b01_100110010010: DATA = 12'b100000000000;
            14'b01_100110010011: DATA = 12'b100000000000;
            14'b01_100110010100: DATA = 12'b100000000000;
            14'b01_100110010101: DATA = 12'b100000000000;
            14'b01_100110010110: DATA = 12'b100000000000;
            14'b01_100110010111: DATA = 12'b100000000000;
            14'b01_100110011000: DATA = 12'b100000000000;
            14'b01_100110011001: DATA = 12'b100000000000;
            14'b01_100110011010: DATA = 12'b100000000000;
            14'b01_100110011011: DATA = 12'b100000000000;
            14'b01_100110011100: DATA = 12'b100000000000;
            14'b01_100110011101: DATA = 12'b100000000000;
            14'b01_100110011110: DATA = 12'b100000000000;
            14'b01_100110011111: DATA = 12'b100000000000;
            14'b01_100110100000: DATA = 12'b100000000000;
            14'b01_100110100001: DATA = 12'b100000000000;
            14'b01_100110100010: DATA = 12'b100000000000;
            14'b01_100110100011: DATA = 12'b100000000000;
            14'b01_100110100100: DATA = 12'b100000000000;
            14'b01_100110100101: DATA = 12'b100000000000;
            14'b01_100110100110: DATA = 12'b100000000000;
            14'b01_100110100111: DATA = 12'b100000000000;
            14'b01_100110101000: DATA = 12'b100000000000;
            14'b01_100110101001: DATA = 12'b100000000000;
            14'b01_100110101010: DATA = 12'b100000000000;
            14'b01_100110101011: DATA = 12'b100000000000;
            14'b01_100110101100: DATA = 12'b100000000000;
            14'b01_100110101101: DATA = 12'b100000000000;
            14'b01_100110101110: DATA = 12'b100000000000;
            14'b01_100110101111: DATA = 12'b100000000000;
            14'b01_100110110000: DATA = 12'b100000000000;
            14'b01_100110110001: DATA = 12'b100000000000;
            14'b01_100110110010: DATA = 12'b100000000000;
            14'b01_100110110011: DATA = 12'b100000000000;
            14'b01_100110110100: DATA = 12'b100000000000;
            14'b01_100110110101: DATA = 12'b100000000000;
            14'b01_100110110110: DATA = 12'b100000000000;
            14'b01_100110110111: DATA = 12'b100000000000;
            14'b01_100110111000: DATA = 12'b100000000000;
            14'b01_100110111001: DATA = 12'b100000000000;
            14'b01_100110111010: DATA = 12'b100000000000;
            14'b01_100110111011: DATA = 12'b100000000000;
            14'b01_100110111100: DATA = 12'b100000000000;
            14'b01_100110111101: DATA = 12'b100000000000;
            14'b01_100110111110: DATA = 12'b100000000000;
            14'b01_100110111111: DATA = 12'b100000000000;
            14'b01_100111000000: DATA = 12'b100000000000;
            14'b01_100111000001: DATA = 12'b100000000000;
            14'b01_100111000010: DATA = 12'b100000000000;
            14'b01_100111000011: DATA = 12'b100000000000;
            14'b01_100111000100: DATA = 12'b100000000000;
            14'b01_100111000101: DATA = 12'b100000000000;
            14'b01_100111000110: DATA = 12'b100000000000;
            14'b01_100111000111: DATA = 12'b100000000000;
            14'b01_100111001000: DATA = 12'b100000000000;
            14'b01_100111001001: DATA = 12'b100000000000;
            14'b01_100111001010: DATA = 12'b100000000000;
            14'b01_100111001011: DATA = 12'b100000000000;
            14'b01_100111001100: DATA = 12'b100000000000;
            14'b01_100111001101: DATA = 12'b100000000000;
            14'b01_100111001110: DATA = 12'b100000000000;
            14'b01_100111001111: DATA = 12'b100000000000;
            14'b01_100111010000: DATA = 12'b100000000000;
            14'b01_100111010001: DATA = 12'b100000000000;
            14'b01_100111010010: DATA = 12'b100000000000;
            14'b01_100111010011: DATA = 12'b100000000000;
            14'b01_100111010100: DATA = 12'b100000000000;
            14'b01_100111010101: DATA = 12'b100000000000;
            14'b01_100111010110: DATA = 12'b100000000000;
            14'b01_100111010111: DATA = 12'b100000000000;
            14'b01_100111011000: DATA = 12'b100000000000;
            14'b01_100111011001: DATA = 12'b100000000000;
            14'b01_100111011010: DATA = 12'b100000000000;
            14'b01_100111011011: DATA = 12'b100000000000;
            14'b01_100111011100: DATA = 12'b100000000000;
            14'b01_100111011101: DATA = 12'b100000000000;
            14'b01_100111011110: DATA = 12'b100000000000;
            14'b01_100111011111: DATA = 12'b100000000000;
            14'b01_100111100000: DATA = 12'b100000000000;
            14'b01_100111100001: DATA = 12'b100000000000;
            14'b01_100111100010: DATA = 12'b100000000000;
            14'b01_100111100011: DATA = 12'b100000000000;
            14'b01_100111100100: DATA = 12'b100000000000;
            14'b01_100111100101: DATA = 12'b100000000000;
            14'b01_100111100110: DATA = 12'b100000000000;
            14'b01_100111100111: DATA = 12'b100000000000;
            14'b01_100111101000: DATA = 12'b100000000000;
            14'b01_100111101001: DATA = 12'b100000000000;
            14'b01_100111101010: DATA = 12'b100000000000;
            14'b01_100111101011: DATA = 12'b100000000000;
            14'b01_100111101100: DATA = 12'b100000000000;
            14'b01_100111101101: DATA = 12'b100000000000;
            14'b01_100111101110: DATA = 12'b100000000000;
            14'b01_100111101111: DATA = 12'b100000000000;
            14'b01_100111110000: DATA = 12'b100000000000;
            14'b01_100111110001: DATA = 12'b100000000000;
            14'b01_100111110010: DATA = 12'b100000000000;
            14'b01_100111110011: DATA = 12'b100000000000;
            14'b01_100111110100: DATA = 12'b100000000000;
            14'b01_100111110101: DATA = 12'b100000000000;
            14'b01_100111110110: DATA = 12'b100000000000;
            14'b01_100111110111: DATA = 12'b100000000000;
            14'b01_100111111000: DATA = 12'b100000000000;
            14'b01_100111111001: DATA = 12'b100000000000;
            14'b01_100111111010: DATA = 12'b100000000000;
            14'b01_100111111011: DATA = 12'b100000000000;
            14'b01_100111111100: DATA = 12'b100000000000;
            14'b01_100111111101: DATA = 12'b100000000000;
            14'b01_100111111110: DATA = 12'b100000000000;
            14'b01_100111111111: DATA = 12'b100000000000;
            14'b01_101000000000: DATA = 12'b100000000000;
            14'b01_101000000001: DATA = 12'b100000000000;
            14'b01_101000000010: DATA = 12'b100000000000;
            14'b01_101000000011: DATA = 12'b100000000000;
            14'b01_101000000100: DATA = 12'b100000000000;
            14'b01_101000000101: DATA = 12'b100000000000;
            14'b01_101000000110: DATA = 12'b100000000000;
            14'b01_101000000111: DATA = 12'b100000000000;
            14'b01_101000001000: DATA = 12'b100000000000;
            14'b01_101000001001: DATA = 12'b100000000000;
            14'b01_101000001010: DATA = 12'b100000000000;
            14'b01_101000001011: DATA = 12'b100000000000;
            14'b01_101000001100: DATA = 12'b100000000000;
            14'b01_101000001101: DATA = 12'b100000000000;
            14'b01_101000001110: DATA = 12'b100000000000;
            14'b01_101000001111: DATA = 12'b100000000000;
            14'b01_101000010000: DATA = 12'b100000000000;
            14'b01_101000010001: DATA = 12'b100000000000;
            14'b01_101000010010: DATA = 12'b100000000000;
            14'b01_101000010011: DATA = 12'b100000000000;
            14'b01_101000010100: DATA = 12'b100000000000;
            14'b01_101000010101: DATA = 12'b100000000000;
            14'b01_101000010110: DATA = 12'b100000000000;
            14'b01_101000010111: DATA = 12'b100000000000;
            14'b01_101000011000: DATA = 12'b100000000000;
            14'b01_101000011001: DATA = 12'b100000000000;
            14'b01_101000011010: DATA = 12'b100000000000;
            14'b01_101000011011: DATA = 12'b100000000000;
            14'b01_101000011100: DATA = 12'b100000000000;
            14'b01_101000011101: DATA = 12'b100000000000;
            14'b01_101000011110: DATA = 12'b100000000000;
            14'b01_101000011111: DATA = 12'b100000000000;
            14'b01_101000100000: DATA = 12'b100000000000;
            14'b01_101000100001: DATA = 12'b100000000000;
            14'b01_101000100010: DATA = 12'b100000000000;
            14'b01_101000100011: DATA = 12'b100000000000;
            14'b01_101000100100: DATA = 12'b100000000000;
            14'b01_101000100101: DATA = 12'b100000000000;
            14'b01_101000100110: DATA = 12'b100000000000;
            14'b01_101000100111: DATA = 12'b100000000000;
            14'b01_101000101000: DATA = 12'b100000000000;
            14'b01_101000101001: DATA = 12'b100000000000;
            14'b01_101000101010: DATA = 12'b100000000000;
            14'b01_101000101011: DATA = 12'b100000000000;
            14'b01_101000101100: DATA = 12'b100000000000;
            14'b01_101000101101: DATA = 12'b100000000000;
            14'b01_101000101110: DATA = 12'b100000000000;
            14'b01_101000101111: DATA = 12'b100000000000;
            14'b01_101000110000: DATA = 12'b100000000000;
            14'b01_101000110001: DATA = 12'b100000000000;
            14'b01_101000110010: DATA = 12'b100000000000;
            14'b01_101000110011: DATA = 12'b100000000000;
            14'b01_101000110100: DATA = 12'b100000000000;
            14'b01_101000110101: DATA = 12'b100000000000;
            14'b01_101000110110: DATA = 12'b100000000000;
            14'b01_101000110111: DATA = 12'b100000000000;
            14'b01_101000111000: DATA = 12'b100000000000;
            14'b01_101000111001: DATA = 12'b100000000000;
            14'b01_101000111010: DATA = 12'b100000000000;
            14'b01_101000111011: DATA = 12'b100000000000;
            14'b01_101000111100: DATA = 12'b100000000000;
            14'b01_101000111101: DATA = 12'b100000000000;
            14'b01_101000111110: DATA = 12'b100000000000;
            14'b01_101000111111: DATA = 12'b100000000000;
            14'b01_101001000000: DATA = 12'b100000000000;
            14'b01_101001000001: DATA = 12'b100000000000;
            14'b01_101001000010: DATA = 12'b100000000000;
            14'b01_101001000011: DATA = 12'b100000000000;
            14'b01_101001000100: DATA = 12'b100000000000;
            14'b01_101001000101: DATA = 12'b100000000000;
            14'b01_101001000110: DATA = 12'b100000000000;
            14'b01_101001000111: DATA = 12'b100000000000;
            14'b01_101001001000: DATA = 12'b100000000000;
            14'b01_101001001001: DATA = 12'b100000000000;
            14'b01_101001001010: DATA = 12'b100000000000;
            14'b01_101001001011: DATA = 12'b100000000000;
            14'b01_101001001100: DATA = 12'b100000000000;
            14'b01_101001001101: DATA = 12'b100000000000;
            14'b01_101001001110: DATA = 12'b100000000000;
            14'b01_101001001111: DATA = 12'b100000000000;
            14'b01_101001010000: DATA = 12'b100000000000;
            14'b01_101001010001: DATA = 12'b100000000000;
            14'b01_101001010010: DATA = 12'b100000000000;
            14'b01_101001010011: DATA = 12'b100000000000;
            14'b01_101001010100: DATA = 12'b100000000000;
            14'b01_101001010101: DATA = 12'b100000000000;
            14'b01_101001010110: DATA = 12'b100000000000;
            14'b01_101001010111: DATA = 12'b100000000000;
            14'b01_101001011000: DATA = 12'b100000000000;
            14'b01_101001011001: DATA = 12'b100000000000;
            14'b01_101001011010: DATA = 12'b100000000000;
            14'b01_101001011011: DATA = 12'b100000000000;
            14'b01_101001011100: DATA = 12'b100000000000;
            14'b01_101001011101: DATA = 12'b100000000000;
            14'b01_101001011110: DATA = 12'b100000000000;
            14'b01_101001011111: DATA = 12'b100000000000;
            14'b01_101001100000: DATA = 12'b100000000000;
            14'b01_101001100001: DATA = 12'b100000000000;
            14'b01_101001100010: DATA = 12'b100000000000;
            14'b01_101001100011: DATA = 12'b100000000000;
            14'b01_101001100100: DATA = 12'b100000000000;
            14'b01_101001100101: DATA = 12'b100000000000;
            14'b01_101001100110: DATA = 12'b100000000000;
            14'b01_101001100111: DATA = 12'b100000000000;
            14'b01_101001101000: DATA = 12'b100000000000;
            14'b01_101001101001: DATA = 12'b100000000000;
            14'b01_101001101010: DATA = 12'b100000000000;
            14'b01_101001101011: DATA = 12'b100000000000;
            14'b01_101001101100: DATA = 12'b100000000000;
            14'b01_101001101101: DATA = 12'b100000000000;
            14'b01_101001101110: DATA = 12'b100000000000;
            14'b01_101001101111: DATA = 12'b100000000000;
            14'b01_101001110000: DATA = 12'b100000000000;
            14'b01_101001110001: DATA = 12'b100000000000;
            14'b01_101001110010: DATA = 12'b100000000000;
            14'b01_101001110011: DATA = 12'b100000000000;
            14'b01_101001110100: DATA = 12'b100000000000;
            14'b01_101001110101: DATA = 12'b100000000000;
            14'b01_101001110110: DATA = 12'b100000000000;
            14'b01_101001110111: DATA = 12'b100000000000;
            14'b01_101001111000: DATA = 12'b100000000000;
            14'b01_101001111001: DATA = 12'b100000000000;
            14'b01_101001111010: DATA = 12'b100000000000;
            14'b01_101001111011: DATA = 12'b100000000000;
            14'b01_101001111100: DATA = 12'b100000000000;
            14'b01_101001111101: DATA = 12'b100000000000;
            14'b01_101001111110: DATA = 12'b100000000000;
            14'b01_101001111111: DATA = 12'b100000000000;
            14'b01_101010000000: DATA = 12'b100000000000;
            14'b01_101010000001: DATA = 12'b100000000000;
            14'b01_101010000010: DATA = 12'b100000000000;
            14'b01_101010000011: DATA = 12'b100000000000;
            14'b01_101010000100: DATA = 12'b100000000000;
            14'b01_101010000101: DATA = 12'b100000000000;
            14'b01_101010000110: DATA = 12'b100000000000;
            14'b01_101010000111: DATA = 12'b100000000000;
            14'b01_101010001000: DATA = 12'b100000000000;
            14'b01_101010001001: DATA = 12'b100000000000;
            14'b01_101010001010: DATA = 12'b100000000000;
            14'b01_101010001011: DATA = 12'b100000000000;
            14'b01_101010001100: DATA = 12'b100000000000;
            14'b01_101010001101: DATA = 12'b100000000000;
            14'b01_101010001110: DATA = 12'b100000000000;
            14'b01_101010001111: DATA = 12'b100000000000;
            14'b01_101010010000: DATA = 12'b100000000000;
            14'b01_101010010001: DATA = 12'b100000000000;
            14'b01_101010010010: DATA = 12'b100000000000;
            14'b01_101010010011: DATA = 12'b100000000000;
            14'b01_101010010100: DATA = 12'b100000000000;
            14'b01_101010010101: DATA = 12'b100000000000;
            14'b01_101010010110: DATA = 12'b100000000000;
            14'b01_101010010111: DATA = 12'b100000000000;
            14'b01_101010011000: DATA = 12'b100000000000;
            14'b01_101010011001: DATA = 12'b100000000000;
            14'b01_101010011010: DATA = 12'b100000000000;
            14'b01_101010011011: DATA = 12'b100000000000;
            14'b01_101010011100: DATA = 12'b100000000000;
            14'b01_101010011101: DATA = 12'b100000000000;
            14'b01_101010011110: DATA = 12'b100000000000;
            14'b01_101010011111: DATA = 12'b100000000000;
            14'b01_101010100000: DATA = 12'b100000000000;
            14'b01_101010100001: DATA = 12'b100000000000;
            14'b01_101010100010: DATA = 12'b100000000000;
            14'b01_101010100011: DATA = 12'b100000000000;
            14'b01_101010100100: DATA = 12'b100000000000;
            14'b01_101010100101: DATA = 12'b100000000000;
            14'b01_101010100110: DATA = 12'b100000000000;
            14'b01_101010100111: DATA = 12'b100000000000;
            14'b01_101010101000: DATA = 12'b100000000000;
            14'b01_101010101001: DATA = 12'b100000000000;
            14'b01_101010101010: DATA = 12'b100000000000;
            14'b01_101010101011: DATA = 12'b100000000000;
            14'b01_101010101100: DATA = 12'b100000000000;
            14'b01_101010101101: DATA = 12'b100000000000;
            14'b01_101010101110: DATA = 12'b100000000000;
            14'b01_101010101111: DATA = 12'b100000000000;
            14'b01_101010110000: DATA = 12'b100000000000;
            14'b01_101010110001: DATA = 12'b100000000000;
            14'b01_101010110010: DATA = 12'b100000000000;
            14'b01_101010110011: DATA = 12'b100000000000;
            14'b01_101010110100: DATA = 12'b100000000000;
            14'b01_101010110101: DATA = 12'b100000000000;
            14'b01_101010110110: DATA = 12'b100000000000;
            14'b01_101010110111: DATA = 12'b100000000000;
            14'b01_101010111000: DATA = 12'b100000000000;
            14'b01_101010111001: DATA = 12'b100000000000;
            14'b01_101010111010: DATA = 12'b100000000000;
            14'b01_101010111011: DATA = 12'b100000000000;
            14'b01_101010111100: DATA = 12'b100000000000;
            14'b01_101010111101: DATA = 12'b100000000000;
            14'b01_101010111110: DATA = 12'b100000000000;
            14'b01_101010111111: DATA = 12'b100000000000;
            14'b01_101011000000: DATA = 12'b100000000000;
            14'b01_101011000001: DATA = 12'b100000000000;
            14'b01_101011000010: DATA = 12'b100000000000;
            14'b01_101011000011: DATA = 12'b100000000000;
            14'b01_101011000100: DATA = 12'b100000000000;
            14'b01_101011000101: DATA = 12'b100000000000;
            14'b01_101011000110: DATA = 12'b100000000000;
            14'b01_101011000111: DATA = 12'b100000000000;
            14'b01_101011001000: DATA = 12'b100000000000;
            14'b01_101011001001: DATA = 12'b100000000000;
            14'b01_101011001010: DATA = 12'b100000000000;
            14'b01_101011001011: DATA = 12'b100000000000;
            14'b01_101011001100: DATA = 12'b100000000000;
            14'b01_101011001101: DATA = 12'b100000000000;
            14'b01_101011001110: DATA = 12'b100000000000;
            14'b01_101011001111: DATA = 12'b100000000000;
            14'b01_101011010000: DATA = 12'b100000000000;
            14'b01_101011010001: DATA = 12'b100000000000;
            14'b01_101011010010: DATA = 12'b100000000000;
            14'b01_101011010011: DATA = 12'b100000000000;
            14'b01_101011010100: DATA = 12'b100000000000;
            14'b01_101011010101: DATA = 12'b100000000000;
            14'b01_101011010110: DATA = 12'b100000000000;
            14'b01_101011010111: DATA = 12'b100000000000;
            14'b01_101011011000: DATA = 12'b100000000000;
            14'b01_101011011001: DATA = 12'b100000000000;
            14'b01_101011011010: DATA = 12'b100000000000;
            14'b01_101011011011: DATA = 12'b100000000000;
            14'b01_101011011100: DATA = 12'b100000000000;
            14'b01_101011011101: DATA = 12'b100000000000;
            14'b01_101011011110: DATA = 12'b100000000000;
            14'b01_101011011111: DATA = 12'b100000000000;
            14'b01_101011100000: DATA = 12'b100000000000;
            14'b01_101011100001: DATA = 12'b100000000000;
            14'b01_101011100010: DATA = 12'b100000000000;
            14'b01_101011100011: DATA = 12'b100000000000;
            14'b01_101011100100: DATA = 12'b100000000000;
            14'b01_101011100101: DATA = 12'b100000000000;
            14'b01_101011100110: DATA = 12'b100000000000;
            14'b01_101011100111: DATA = 12'b100000000000;
            14'b01_101011101000: DATA = 12'b100000000000;
            14'b01_101011101001: DATA = 12'b100000000000;
            14'b01_101011101010: DATA = 12'b100000000000;
            14'b01_101011101011: DATA = 12'b100000000000;
            14'b01_101011101100: DATA = 12'b100000000000;
            14'b01_101011101101: DATA = 12'b100000000000;
            14'b01_101011101110: DATA = 12'b100000000000;
            14'b01_101011101111: DATA = 12'b100000000000;
            14'b01_101011110000: DATA = 12'b100000000000;
            14'b01_101011110001: DATA = 12'b100000000000;
            14'b01_101011110010: DATA = 12'b100000000000;
            14'b01_101011110011: DATA = 12'b100000000000;
            14'b01_101011110100: DATA = 12'b100000000000;
            14'b01_101011110101: DATA = 12'b100000000000;
            14'b01_101011110110: DATA = 12'b100000000000;
            14'b01_101011110111: DATA = 12'b100000000000;
            14'b01_101011111000: DATA = 12'b100000000000;
            14'b01_101011111001: DATA = 12'b100000000000;
            14'b01_101011111010: DATA = 12'b100000000000;
            14'b01_101011111011: DATA = 12'b100000000000;
            14'b01_101011111100: DATA = 12'b100000000000;
            14'b01_101011111101: DATA = 12'b100000000000;
            14'b01_101011111110: DATA = 12'b100000000000;
            14'b01_101011111111: DATA = 12'b100000000000;
            14'b01_101100000000: DATA = 12'b100000000000;
            14'b01_101100000001: DATA = 12'b100000000000;
            14'b01_101100000010: DATA = 12'b100000000000;
            14'b01_101100000011: DATA = 12'b100000000000;
            14'b01_101100000100: DATA = 12'b100000000000;
            14'b01_101100000101: DATA = 12'b100000000000;
            14'b01_101100000110: DATA = 12'b100000000000;
            14'b01_101100000111: DATA = 12'b100000000000;
            14'b01_101100001000: DATA = 12'b100000000000;
            14'b01_101100001001: DATA = 12'b100000000000;
            14'b01_101100001010: DATA = 12'b100000000000;
            14'b01_101100001011: DATA = 12'b100000000000;
            14'b01_101100001100: DATA = 12'b100000000000;
            14'b01_101100001101: DATA = 12'b100000000000;
            14'b01_101100001110: DATA = 12'b100000000000;
            14'b01_101100001111: DATA = 12'b100000000000;
            14'b01_101100010000: DATA = 12'b100000000000;
            14'b01_101100010001: DATA = 12'b100000000000;
            14'b01_101100010010: DATA = 12'b100000000000;
            14'b01_101100010011: DATA = 12'b100000000000;
            14'b01_101100010100: DATA = 12'b100000000000;
            14'b01_101100010101: DATA = 12'b100000000000;
            14'b01_101100010110: DATA = 12'b100000000000;
            14'b01_101100010111: DATA = 12'b100000000000;
            14'b01_101100011000: DATA = 12'b100000000000;
            14'b01_101100011001: DATA = 12'b100000000000;
            14'b01_101100011010: DATA = 12'b100000000000;
            14'b01_101100011011: DATA = 12'b100000000000;
            14'b01_101100011100: DATA = 12'b100000000000;
            14'b01_101100011101: DATA = 12'b100000000000;
            14'b01_101100011110: DATA = 12'b100000000000;
            14'b01_101100011111: DATA = 12'b100000000000;
            14'b01_101100100000: DATA = 12'b100000000000;
            14'b01_101100100001: DATA = 12'b100000000000;
            14'b01_101100100010: DATA = 12'b100000000000;
            14'b01_101100100011: DATA = 12'b100000000000;
            14'b01_101100100100: DATA = 12'b100000000000;
            14'b01_101100100101: DATA = 12'b100000000000;
            14'b01_101100100110: DATA = 12'b100000000000;
            14'b01_101100100111: DATA = 12'b100000000000;
            14'b01_101100101000: DATA = 12'b100000000000;
            14'b01_101100101001: DATA = 12'b100000000000;
            14'b01_101100101010: DATA = 12'b100000000000;
            14'b01_101100101011: DATA = 12'b100000000000;
            14'b01_101100101100: DATA = 12'b100000000000;
            14'b01_101100101101: DATA = 12'b100000000000;
            14'b01_101100101110: DATA = 12'b100000000000;
            14'b01_101100101111: DATA = 12'b100000000000;
            14'b01_101100110000: DATA = 12'b100000000000;
            14'b01_101100110001: DATA = 12'b100000000000;
            14'b01_101100110010: DATA = 12'b100000000000;
            14'b01_101100110011: DATA = 12'b100000000000;
            14'b01_101100110100: DATA = 12'b100000000000;
            14'b01_101100110101: DATA = 12'b100000000000;
            14'b01_101100110110: DATA = 12'b100000000000;
            14'b01_101100110111: DATA = 12'b100000000000;
            14'b01_101100111000: DATA = 12'b100000000000;
            14'b01_101100111001: DATA = 12'b100000000000;
            14'b01_101100111010: DATA = 12'b100000000000;
            14'b01_101100111011: DATA = 12'b100000000000;
            14'b01_101100111100: DATA = 12'b100000000000;
            14'b01_101100111101: DATA = 12'b100000000000;
            14'b01_101100111110: DATA = 12'b100000000000;
            14'b01_101100111111: DATA = 12'b100000000000;
            14'b01_101101000000: DATA = 12'b100000000000;
            14'b01_101101000001: DATA = 12'b100000000000;
            14'b01_101101000010: DATA = 12'b100000000000;
            14'b01_101101000011: DATA = 12'b100000000000;
            14'b01_101101000100: DATA = 12'b100000000000;
            14'b01_101101000101: DATA = 12'b100000000000;
            14'b01_101101000110: DATA = 12'b100000000000;
            14'b01_101101000111: DATA = 12'b100000000000;
            14'b01_101101001000: DATA = 12'b100000000000;
            14'b01_101101001001: DATA = 12'b100000000000;
            14'b01_101101001010: DATA = 12'b100000000000;
            14'b01_101101001011: DATA = 12'b100000000000;
            14'b01_101101001100: DATA = 12'b100000000000;
            14'b01_101101001101: DATA = 12'b100000000000;
            14'b01_101101001110: DATA = 12'b100000000000;
            14'b01_101101001111: DATA = 12'b100000000000;
            14'b01_101101010000: DATA = 12'b100000000000;
            14'b01_101101010001: DATA = 12'b100000000000;
            14'b01_101101010010: DATA = 12'b100000000000;
            14'b01_101101010011: DATA = 12'b100000000000;
            14'b01_101101010100: DATA = 12'b100000000000;
            14'b01_101101010101: DATA = 12'b100000000000;
            14'b01_101101010110: DATA = 12'b100000000000;
            14'b01_101101010111: DATA = 12'b100000000000;
            14'b01_101101011000: DATA = 12'b100000000000;
            14'b01_101101011001: DATA = 12'b100000000000;
            14'b01_101101011010: DATA = 12'b100000000000;
            14'b01_101101011011: DATA = 12'b100000000000;
            14'b01_101101011100: DATA = 12'b100000000000;
            14'b01_101101011101: DATA = 12'b100000000000;
            14'b01_101101011110: DATA = 12'b100000000000;
            14'b01_101101011111: DATA = 12'b100000000000;
            14'b01_101101100000: DATA = 12'b100000000000;
            14'b01_101101100001: DATA = 12'b100000000000;
            14'b01_101101100010: DATA = 12'b100000000000;
            14'b01_101101100011: DATA = 12'b100000000000;
            14'b01_101101100100: DATA = 12'b100000000000;
            14'b01_101101100101: DATA = 12'b100000000000;
            14'b01_101101100110: DATA = 12'b100000000000;
            14'b01_101101100111: DATA = 12'b100000000000;
            14'b01_101101101000: DATA = 12'b100000000000;
            14'b01_101101101001: DATA = 12'b100000000000;
            14'b01_101101101010: DATA = 12'b100000000000;
            14'b01_101101101011: DATA = 12'b100000000000;
            14'b01_101101101100: DATA = 12'b100000000000;
            14'b01_101101101101: DATA = 12'b100000000000;
            14'b01_101101101110: DATA = 12'b100000000000;
            14'b01_101101101111: DATA = 12'b100000000000;
            14'b01_101101110000: DATA = 12'b100000000000;
            14'b01_101101110001: DATA = 12'b100000000000;
            14'b01_101101110010: DATA = 12'b100000000000;
            14'b01_101101110011: DATA = 12'b100000000000;
            14'b01_101101110100: DATA = 12'b100000000000;
            14'b01_101101110101: DATA = 12'b100000000000;
            14'b01_101101110110: DATA = 12'b100000000000;
            14'b01_101101110111: DATA = 12'b100000000000;
            14'b01_101101111000: DATA = 12'b100000000000;
            14'b01_101101111001: DATA = 12'b100000000000;
            14'b01_101101111010: DATA = 12'b100000000000;
            14'b01_101101111011: DATA = 12'b100000000000;
            14'b01_101101111100: DATA = 12'b100000000000;
            14'b01_101101111101: DATA = 12'b100000000000;
            14'b01_101101111110: DATA = 12'b100000000000;
            14'b01_101101111111: DATA = 12'b100000000000;
            14'b01_101110000000: DATA = 12'b100000000000;
            14'b01_101110000001: DATA = 12'b100000000000;
            14'b01_101110000010: DATA = 12'b100000000000;
            14'b01_101110000011: DATA = 12'b100000000000;
            14'b01_101110000100: DATA = 12'b100000000000;
            14'b01_101110000101: DATA = 12'b100000000000;
            14'b01_101110000110: DATA = 12'b100000000000;
            14'b01_101110000111: DATA = 12'b100000000000;
            14'b01_101110001000: DATA = 12'b100000000000;
            14'b01_101110001001: DATA = 12'b100000000000;
            14'b01_101110001010: DATA = 12'b100000000000;
            14'b01_101110001011: DATA = 12'b100000000000;
            14'b01_101110001100: DATA = 12'b100000000000;
            14'b01_101110001101: DATA = 12'b100000000000;
            14'b01_101110001110: DATA = 12'b100000000000;
            14'b01_101110001111: DATA = 12'b100000000000;
            14'b01_101110010000: DATA = 12'b100000000000;
            14'b01_101110010001: DATA = 12'b100000000000;
            14'b01_101110010010: DATA = 12'b100000000000;
            14'b01_101110010011: DATA = 12'b100000000000;
            14'b01_101110010100: DATA = 12'b100000000000;
            14'b01_101110010101: DATA = 12'b100000000000;
            14'b01_101110010110: DATA = 12'b100000000000;
            14'b01_101110010111: DATA = 12'b100000000000;
            14'b01_101110011000: DATA = 12'b100000000000;
            14'b01_101110011001: DATA = 12'b100000000000;
            14'b01_101110011010: DATA = 12'b100000000000;
            14'b01_101110011011: DATA = 12'b100000000000;
            14'b01_101110011100: DATA = 12'b100000000000;
            14'b01_101110011101: DATA = 12'b100000000000;
            14'b01_101110011110: DATA = 12'b100000000000;
            14'b01_101110011111: DATA = 12'b100000000000;
            14'b01_101110100000: DATA = 12'b100000000000;
            14'b01_101110100001: DATA = 12'b100000000000;
            14'b01_101110100010: DATA = 12'b100000000000;
            14'b01_101110100011: DATA = 12'b100000000000;
            14'b01_101110100100: DATA = 12'b100000000000;
            14'b01_101110100101: DATA = 12'b100000000000;
            14'b01_101110100110: DATA = 12'b100000000000;
            14'b01_101110100111: DATA = 12'b100000000000;
            14'b01_101110101000: DATA = 12'b100000000000;
            14'b01_101110101001: DATA = 12'b100000000000;
            14'b01_101110101010: DATA = 12'b100000000000;
            14'b01_101110101011: DATA = 12'b100000000000;
            14'b01_101110101100: DATA = 12'b100000000000;
            14'b01_101110101101: DATA = 12'b100000000000;
            14'b01_101110101110: DATA = 12'b100000000000;
            14'b01_101110101111: DATA = 12'b100000000000;
            14'b01_101110110000: DATA = 12'b100000000000;
            14'b01_101110110001: DATA = 12'b100000000000;
            14'b01_101110110010: DATA = 12'b100000000000;
            14'b01_101110110011: DATA = 12'b100000000000;
            14'b01_101110110100: DATA = 12'b100000000000;
            14'b01_101110110101: DATA = 12'b100000000000;
            14'b01_101110110110: DATA = 12'b100000000000;
            14'b01_101110110111: DATA = 12'b100000000000;
            14'b01_101110111000: DATA = 12'b100000000000;
            14'b01_101110111001: DATA = 12'b100000000000;
            14'b01_101110111010: DATA = 12'b100000000000;
            14'b01_101110111011: DATA = 12'b100000000000;
            14'b01_101110111100: DATA = 12'b100000000000;
            14'b01_101110111101: DATA = 12'b100000000000;
            14'b01_101110111110: DATA = 12'b100000000000;
            14'b01_101110111111: DATA = 12'b100000000000;
            14'b01_101111000000: DATA = 12'b100000000000;
            14'b01_101111000001: DATA = 12'b100000000000;
            14'b01_101111000010: DATA = 12'b100000000000;
            14'b01_101111000011: DATA = 12'b100000000000;
            14'b01_101111000100: DATA = 12'b100000000000;
            14'b01_101111000101: DATA = 12'b100000000000;
            14'b01_101111000110: DATA = 12'b100000000000;
            14'b01_101111000111: DATA = 12'b100000000000;
            14'b01_101111001000: DATA = 12'b100000000000;
            14'b01_101111001001: DATA = 12'b100000000000;
            14'b01_101111001010: DATA = 12'b100000000000;
            14'b01_101111001011: DATA = 12'b100000000000;
            14'b01_101111001100: DATA = 12'b100000000000;
            14'b01_101111001101: DATA = 12'b100000000000;
            14'b01_101111001110: DATA = 12'b100000000000;
            14'b01_101111001111: DATA = 12'b100000000000;
            14'b01_101111010000: DATA = 12'b100000000000;
            14'b01_101111010001: DATA = 12'b100000000000;
            14'b01_101111010010: DATA = 12'b100000000000;
            14'b01_101111010011: DATA = 12'b100000000000;
            14'b01_101111010100: DATA = 12'b100000000000;
            14'b01_101111010101: DATA = 12'b100000000000;
            14'b01_101111010110: DATA = 12'b100000000000;
            14'b01_101111010111: DATA = 12'b100000000000;
            14'b01_101111011000: DATA = 12'b100000000000;
            14'b01_101111011001: DATA = 12'b100000000000;
            14'b01_101111011010: DATA = 12'b100000000000;
            14'b01_101111011011: DATA = 12'b100000000000;
            14'b01_101111011100: DATA = 12'b100000000000;
            14'b01_101111011101: DATA = 12'b100000000000;
            14'b01_101111011110: DATA = 12'b100000000000;
            14'b01_101111011111: DATA = 12'b100000000000;
            14'b01_101111100000: DATA = 12'b100000000000;
            14'b01_101111100001: DATA = 12'b100000000000;
            14'b01_101111100010: DATA = 12'b100000000000;
            14'b01_101111100011: DATA = 12'b100000000000;
            14'b01_101111100100: DATA = 12'b100000000000;
            14'b01_101111100101: DATA = 12'b100000000000;
            14'b01_101111100110: DATA = 12'b100000000000;
            14'b01_101111100111: DATA = 12'b100000000000;
            14'b01_101111101000: DATA = 12'b100000000000;
            14'b01_101111101001: DATA = 12'b100000000000;
            14'b01_101111101010: DATA = 12'b100000000000;
            14'b01_101111101011: DATA = 12'b100000000000;
            14'b01_101111101100: DATA = 12'b100000000000;
            14'b01_101111101101: DATA = 12'b100000000000;
            14'b01_101111101110: DATA = 12'b100000000000;
            14'b01_101111101111: DATA = 12'b100000000000;
            14'b01_101111110000: DATA = 12'b100000000000;
            14'b01_101111110001: DATA = 12'b100000000000;
            14'b01_101111110010: DATA = 12'b100000000000;
            14'b01_101111110011: DATA = 12'b100000000000;
            14'b01_101111110100: DATA = 12'b100000000000;
            14'b01_101111110101: DATA = 12'b100000000000;
            14'b01_101111110110: DATA = 12'b100000000000;
            14'b01_101111110111: DATA = 12'b100000000000;
            14'b01_101111111000: DATA = 12'b100000000000;
            14'b01_101111111001: DATA = 12'b100000000000;
            14'b01_101111111010: DATA = 12'b100000000000;
            14'b01_101111111011: DATA = 12'b100000000000;
            14'b01_101111111100: DATA = 12'b100000000000;
            14'b01_101111111101: DATA = 12'b100000000000;
            14'b01_101111111110: DATA = 12'b100000000000;
            14'b01_101111111111: DATA = 12'b100000000000;
            14'b01_110000000000: DATA = 12'b100000000000;
            14'b01_110000000001: DATA = 12'b100000000000;
            14'b01_110000000010: DATA = 12'b100000000000;
            14'b01_110000000011: DATA = 12'b100000000000;
            14'b01_110000000100: DATA = 12'b100000000000;
            14'b01_110000000101: DATA = 12'b100000000000;
            14'b01_110000000110: DATA = 12'b100000000000;
            14'b01_110000000111: DATA = 12'b100000000000;
            14'b01_110000001000: DATA = 12'b100000000000;
            14'b01_110000001001: DATA = 12'b100000000000;
            14'b01_110000001010: DATA = 12'b100000000000;
            14'b01_110000001011: DATA = 12'b100000000000;
            14'b01_110000001100: DATA = 12'b100000000000;
            14'b01_110000001101: DATA = 12'b100000000000;
            14'b01_110000001110: DATA = 12'b100000000000;
            14'b01_110000001111: DATA = 12'b100000000000;
            14'b01_110000010000: DATA = 12'b100000000000;
            14'b01_110000010001: DATA = 12'b100000000000;
            14'b01_110000010010: DATA = 12'b100000000000;
            14'b01_110000010011: DATA = 12'b100000000000;
            14'b01_110000010100: DATA = 12'b100000000000;
            14'b01_110000010101: DATA = 12'b100000000000;
            14'b01_110000010110: DATA = 12'b100000000000;
            14'b01_110000010111: DATA = 12'b100000000000;
            14'b01_110000011000: DATA = 12'b100000000000;
            14'b01_110000011001: DATA = 12'b100000000000;
            14'b01_110000011010: DATA = 12'b100000000000;
            14'b01_110000011011: DATA = 12'b100000000000;
            14'b01_110000011100: DATA = 12'b100000000000;
            14'b01_110000011101: DATA = 12'b100000000000;
            14'b01_110000011110: DATA = 12'b100000000000;
            14'b01_110000011111: DATA = 12'b100000000000;
            14'b01_110000100000: DATA = 12'b100000000000;
            14'b01_110000100001: DATA = 12'b100000000000;
            14'b01_110000100010: DATA = 12'b100000000000;
            14'b01_110000100011: DATA = 12'b100000000000;
            14'b01_110000100100: DATA = 12'b100000000000;
            14'b01_110000100101: DATA = 12'b100000000000;
            14'b01_110000100110: DATA = 12'b100000000000;
            14'b01_110000100111: DATA = 12'b100000000000;
            14'b01_110000101000: DATA = 12'b100000000000;
            14'b01_110000101001: DATA = 12'b100000000000;
            14'b01_110000101010: DATA = 12'b100000000000;
            14'b01_110000101011: DATA = 12'b100000000000;
            14'b01_110000101100: DATA = 12'b100000000000;
            14'b01_110000101101: DATA = 12'b100000000000;
            14'b01_110000101110: DATA = 12'b100000000000;
            14'b01_110000101111: DATA = 12'b100000000000;
            14'b01_110000110000: DATA = 12'b100000000000;
            14'b01_110000110001: DATA = 12'b100000000000;
            14'b01_110000110010: DATA = 12'b100000000000;
            14'b01_110000110011: DATA = 12'b100000000000;
            14'b01_110000110100: DATA = 12'b100000000000;
            14'b01_110000110101: DATA = 12'b100000000000;
            14'b01_110000110110: DATA = 12'b100000000000;
            14'b01_110000110111: DATA = 12'b100000000000;
            14'b01_110000111000: DATA = 12'b100000000000;
            14'b01_110000111001: DATA = 12'b100000000000;
            14'b01_110000111010: DATA = 12'b100000000000;
            14'b01_110000111011: DATA = 12'b100000000000;
            14'b01_110000111100: DATA = 12'b100000000000;
            14'b01_110000111101: DATA = 12'b100000000000;
            14'b01_110000111110: DATA = 12'b100000000000;
            14'b01_110000111111: DATA = 12'b100000000000;
            14'b01_110001000000: DATA = 12'b100000000000;
            14'b01_110001000001: DATA = 12'b100000000000;
            14'b01_110001000010: DATA = 12'b100000000000;
            14'b01_110001000011: DATA = 12'b100000000000;
            14'b01_110001000100: DATA = 12'b100000000000;
            14'b01_110001000101: DATA = 12'b100000000000;
            14'b01_110001000110: DATA = 12'b100000000000;
            14'b01_110001000111: DATA = 12'b100000000000;
            14'b01_110001001000: DATA = 12'b100000000000;
            14'b01_110001001001: DATA = 12'b100000000000;
            14'b01_110001001010: DATA = 12'b100000000000;
            14'b01_110001001011: DATA = 12'b100000000000;
            14'b01_110001001100: DATA = 12'b100000000000;
            14'b01_110001001101: DATA = 12'b100000000000;
            14'b01_110001001110: DATA = 12'b100000000000;
            14'b01_110001001111: DATA = 12'b100000000000;
            14'b01_110001010000: DATA = 12'b100000000000;
            14'b01_110001010001: DATA = 12'b100000000000;
            14'b01_110001010010: DATA = 12'b100000000000;
            14'b01_110001010011: DATA = 12'b100000000000;
            14'b01_110001010100: DATA = 12'b100000000000;
            14'b01_110001010101: DATA = 12'b100000000000;
            14'b01_110001010110: DATA = 12'b100000000000;
            14'b01_110001010111: DATA = 12'b100000000000;
            14'b01_110001011000: DATA = 12'b100000000000;
            14'b01_110001011001: DATA = 12'b100000000000;
            14'b01_110001011010: DATA = 12'b100000000000;
            14'b01_110001011011: DATA = 12'b100000000000;
            14'b01_110001011100: DATA = 12'b100000000000;
            14'b01_110001011101: DATA = 12'b100000000000;
            14'b01_110001011110: DATA = 12'b100000000000;
            14'b01_110001011111: DATA = 12'b100000000000;
            14'b01_110001100000: DATA = 12'b100000000000;
            14'b01_110001100001: DATA = 12'b100000000000;
            14'b01_110001100010: DATA = 12'b100000000000;
            14'b01_110001100011: DATA = 12'b100000000000;
            14'b01_110001100100: DATA = 12'b100000000000;
            14'b01_110001100101: DATA = 12'b100000000000;
            14'b01_110001100110: DATA = 12'b100000000000;
            14'b01_110001100111: DATA = 12'b100000000000;
            14'b01_110001101000: DATA = 12'b100000000000;
            14'b01_110001101001: DATA = 12'b100000000000;
            14'b01_110001101010: DATA = 12'b100000000000;
            14'b01_110001101011: DATA = 12'b100000000000;
            14'b01_110001101100: DATA = 12'b100000000000;
            14'b01_110001101101: DATA = 12'b100000000000;
            14'b01_110001101110: DATA = 12'b100000000000;
            14'b01_110001101111: DATA = 12'b100000000000;
            14'b01_110001110000: DATA = 12'b100000000000;
            14'b01_110001110001: DATA = 12'b100000000000;
            14'b01_110001110010: DATA = 12'b100000000000;
            14'b01_110001110011: DATA = 12'b100000000000;
            14'b01_110001110100: DATA = 12'b100000000000;
            14'b01_110001110101: DATA = 12'b100000000000;
            14'b01_110001110110: DATA = 12'b100000000000;
            14'b01_110001110111: DATA = 12'b100000000000;
            14'b01_110001111000: DATA = 12'b100000000000;
            14'b01_110001111001: DATA = 12'b100000000000;
            14'b01_110001111010: DATA = 12'b100000000000;
            14'b01_110001111011: DATA = 12'b100000000000;
            14'b01_110001111100: DATA = 12'b100000000000;
            14'b01_110001111101: DATA = 12'b100000000000;
            14'b01_110001111110: DATA = 12'b100000000000;
            14'b01_110001111111: DATA = 12'b100000000000;
            14'b01_110010000000: DATA = 12'b100000000000;
            14'b01_110010000001: DATA = 12'b100000000000;
            14'b01_110010000010: DATA = 12'b100000000000;
            14'b01_110010000011: DATA = 12'b100000000000;
            14'b01_110010000100: DATA = 12'b100000000000;
            14'b01_110010000101: DATA = 12'b100000000000;
            14'b01_110010000110: DATA = 12'b100000000000;
            14'b01_110010000111: DATA = 12'b100000000000;
            14'b01_110010001000: DATA = 12'b100000000000;
            14'b01_110010001001: DATA = 12'b100000000000;
            14'b01_110010001010: DATA = 12'b100000000000;
            14'b01_110010001011: DATA = 12'b100000000000;
            14'b01_110010001100: DATA = 12'b100000000000;
            14'b01_110010001101: DATA = 12'b100000000000;
            14'b01_110010001110: DATA = 12'b100000000000;
            14'b01_110010001111: DATA = 12'b100000000000;
            14'b01_110010010000: DATA = 12'b100000000000;
            14'b01_110010010001: DATA = 12'b100000000000;
            14'b01_110010010010: DATA = 12'b100000000000;
            14'b01_110010010011: DATA = 12'b100000000000;
            14'b01_110010010100: DATA = 12'b100000000000;
            14'b01_110010010101: DATA = 12'b100000000000;
            14'b01_110010010110: DATA = 12'b100000000000;
            14'b01_110010010111: DATA = 12'b100000000000;
            14'b01_110010011000: DATA = 12'b100000000000;
            14'b01_110010011001: DATA = 12'b100000000000;
            14'b01_110010011010: DATA = 12'b100000000000;
            14'b01_110010011011: DATA = 12'b100000000000;
            14'b01_110010011100: DATA = 12'b100000000000;
            14'b01_110010011101: DATA = 12'b100000000000;
            14'b01_110010011110: DATA = 12'b100000000000;
            14'b01_110010011111: DATA = 12'b100000000000;
            14'b01_110010100000: DATA = 12'b100000000000;
            14'b01_110010100001: DATA = 12'b100000000000;
            14'b01_110010100010: DATA = 12'b100000000000;
            14'b01_110010100011: DATA = 12'b100000000000;
            14'b01_110010100100: DATA = 12'b100000000000;
            14'b01_110010100101: DATA = 12'b100000000000;
            14'b01_110010100110: DATA = 12'b100000000000;
            14'b01_110010100111: DATA = 12'b100000000000;
            14'b01_110010101000: DATA = 12'b100000000000;
            14'b01_110010101001: DATA = 12'b100000000000;
            14'b01_110010101010: DATA = 12'b100000000000;
            14'b01_110010101011: DATA = 12'b100000000000;
            14'b01_110010101100: DATA = 12'b100000000000;
            14'b01_110010101101: DATA = 12'b100000000000;
            14'b01_110010101110: DATA = 12'b100000000000;
            14'b01_110010101111: DATA = 12'b100000000000;
            14'b01_110010110000: DATA = 12'b100000000000;
            14'b01_110010110001: DATA = 12'b100000000000;
            14'b01_110010110010: DATA = 12'b100000000000;
            14'b01_110010110011: DATA = 12'b100000000000;
            14'b01_110010110100: DATA = 12'b100000000000;
            14'b01_110010110101: DATA = 12'b100000000000;
            14'b01_110010110110: DATA = 12'b100000000000;
            14'b01_110010110111: DATA = 12'b100000000000;
            14'b01_110010111000: DATA = 12'b100000000000;
            14'b01_110010111001: DATA = 12'b100000000000;
            14'b01_110010111010: DATA = 12'b100000000000;
            14'b01_110010111011: DATA = 12'b100000000000;
            14'b01_110010111100: DATA = 12'b100000000000;
            14'b01_110010111101: DATA = 12'b100000000000;
            14'b01_110010111110: DATA = 12'b100000000000;
            14'b01_110010111111: DATA = 12'b100000000000;
            14'b01_110011000000: DATA = 12'b100000000000;
            14'b01_110011000001: DATA = 12'b100000000000;
            14'b01_110011000010: DATA = 12'b100000000000;
            14'b01_110011000011: DATA = 12'b100000000000;
            14'b01_110011000100: DATA = 12'b100000000000;
            14'b01_110011000101: DATA = 12'b100000000000;
            14'b01_110011000110: DATA = 12'b100000000000;
            14'b01_110011000111: DATA = 12'b100000000000;
            14'b01_110011001000: DATA = 12'b100000000000;
            14'b01_110011001001: DATA = 12'b100000000000;
            14'b01_110011001010: DATA = 12'b100000000000;
            14'b01_110011001011: DATA = 12'b100000000000;
            14'b01_110011001100: DATA = 12'b100000000000;
            14'b01_110011001101: DATA = 12'b100000000000;
            14'b01_110011001110: DATA = 12'b100000000000;
            14'b01_110011001111: DATA = 12'b100000000000;
            14'b01_110011010000: DATA = 12'b100000000000;
            14'b01_110011010001: DATA = 12'b100000000000;
            14'b01_110011010010: DATA = 12'b100000000000;
            14'b01_110011010011: DATA = 12'b100000000000;
            14'b01_110011010100: DATA = 12'b100000000000;
            14'b01_110011010101: DATA = 12'b100000000000;
            14'b01_110011010110: DATA = 12'b100000000000;
            14'b01_110011010111: DATA = 12'b100000000000;
            14'b01_110011011000: DATA = 12'b100000000000;
            14'b01_110011011001: DATA = 12'b100000000000;
            14'b01_110011011010: DATA = 12'b100000000000;
            14'b01_110011011011: DATA = 12'b100000000000;
            14'b01_110011011100: DATA = 12'b100000000000;
            14'b01_110011011101: DATA = 12'b100000000000;
            14'b01_110011011110: DATA = 12'b100000000000;
            14'b01_110011011111: DATA = 12'b100000000000;
            14'b01_110011100000: DATA = 12'b100000000000;
            14'b01_110011100001: DATA = 12'b100000000000;
            14'b01_110011100010: DATA = 12'b100000000000;
            14'b01_110011100011: DATA = 12'b100000000000;
            14'b01_110011100100: DATA = 12'b100000000000;
            14'b01_110011100101: DATA = 12'b100000000000;
            14'b01_110011100110: DATA = 12'b100000000000;
            14'b01_110011100111: DATA = 12'b100000000000;
            14'b01_110011101000: DATA = 12'b100000000000;
            14'b01_110011101001: DATA = 12'b100000000000;
            14'b01_110011101010: DATA = 12'b100000000000;
            14'b01_110011101011: DATA = 12'b100000000000;
            14'b01_110011101100: DATA = 12'b100000000000;
            14'b01_110011101101: DATA = 12'b100000000000;
            14'b01_110011101110: DATA = 12'b100000000000;
            14'b01_110011101111: DATA = 12'b100000000000;
            14'b01_110011110000: DATA = 12'b100000000000;
            14'b01_110011110001: DATA = 12'b100000000000;
            14'b01_110011110010: DATA = 12'b100000000000;
            14'b01_110011110011: DATA = 12'b100000000000;
            14'b01_110011110100: DATA = 12'b100000000000;
            14'b01_110011110101: DATA = 12'b100000000000;
            14'b01_110011110110: DATA = 12'b100000000000;
            14'b01_110011110111: DATA = 12'b100000000000;
            14'b01_110011111000: DATA = 12'b100000000000;
            14'b01_110011111001: DATA = 12'b100000000000;
            14'b01_110011111010: DATA = 12'b100000000000;
            14'b01_110011111011: DATA = 12'b100000000000;
            14'b01_110011111100: DATA = 12'b100000000000;
            14'b01_110011111101: DATA = 12'b100000000000;
            14'b01_110011111110: DATA = 12'b100000000000;
            14'b01_110011111111: DATA = 12'b100000000000;
            14'b01_110100000000: DATA = 12'b100000000000;
            14'b01_110100000001: DATA = 12'b100000000000;
            14'b01_110100000010: DATA = 12'b100000000000;
            14'b01_110100000011: DATA = 12'b100000000000;
            14'b01_110100000100: DATA = 12'b100000000000;
            14'b01_110100000101: DATA = 12'b100000000000;
            14'b01_110100000110: DATA = 12'b100000000000;
            14'b01_110100000111: DATA = 12'b100000000000;
            14'b01_110100001000: DATA = 12'b100000000000;
            14'b01_110100001001: DATA = 12'b100000000000;
            14'b01_110100001010: DATA = 12'b100000000000;
            14'b01_110100001011: DATA = 12'b100000000000;
            14'b01_110100001100: DATA = 12'b100000000000;
            14'b01_110100001101: DATA = 12'b100000000000;
            14'b01_110100001110: DATA = 12'b100000000000;
            14'b01_110100001111: DATA = 12'b100000000000;
            14'b01_110100010000: DATA = 12'b100000000000;
            14'b01_110100010001: DATA = 12'b100000000000;
            14'b01_110100010010: DATA = 12'b100000000000;
            14'b01_110100010011: DATA = 12'b100000000000;
            14'b01_110100010100: DATA = 12'b100000000000;
            14'b01_110100010101: DATA = 12'b100000000000;
            14'b01_110100010110: DATA = 12'b100000000000;
            14'b01_110100010111: DATA = 12'b100000000000;
            14'b01_110100011000: DATA = 12'b100000000000;
            14'b01_110100011001: DATA = 12'b100000000000;
            14'b01_110100011010: DATA = 12'b100000000000;
            14'b01_110100011011: DATA = 12'b100000000000;
            14'b01_110100011100: DATA = 12'b100000000000;
            14'b01_110100011101: DATA = 12'b100000000000;
            14'b01_110100011110: DATA = 12'b100000000000;
            14'b01_110100011111: DATA = 12'b100000000000;
            14'b01_110100100000: DATA = 12'b100000000000;
            14'b01_110100100001: DATA = 12'b100000000000;
            14'b01_110100100010: DATA = 12'b100000000000;
            14'b01_110100100011: DATA = 12'b100000000000;
            14'b01_110100100100: DATA = 12'b100000000000;
            14'b01_110100100101: DATA = 12'b100000000000;
            14'b01_110100100110: DATA = 12'b100000000000;
            14'b01_110100100111: DATA = 12'b100000000000;
            14'b01_110100101000: DATA = 12'b100000000000;
            14'b01_110100101001: DATA = 12'b100000000000;
            14'b01_110100101010: DATA = 12'b100000000000;
            14'b01_110100101011: DATA = 12'b100000000000;
            14'b01_110100101100: DATA = 12'b100000000000;
            14'b01_110100101101: DATA = 12'b100000000000;
            14'b01_110100101110: DATA = 12'b100000000000;
            14'b01_110100101111: DATA = 12'b100000000000;
            14'b01_110100110000: DATA = 12'b100000000000;
            14'b01_110100110001: DATA = 12'b100000000000;
            14'b01_110100110010: DATA = 12'b100000000000;
            14'b01_110100110011: DATA = 12'b100000000000;
            14'b01_110100110100: DATA = 12'b100000000000;
            14'b01_110100110101: DATA = 12'b100000000000;
            14'b01_110100110110: DATA = 12'b100000000000;
            14'b01_110100110111: DATA = 12'b100000000000;
            14'b01_110100111000: DATA = 12'b100000000000;
            14'b01_110100111001: DATA = 12'b100000000000;
            14'b01_110100111010: DATA = 12'b100000000000;
            14'b01_110100111011: DATA = 12'b100000000000;
            14'b01_110100111100: DATA = 12'b100000000000;
            14'b01_110100111101: DATA = 12'b100000000000;
            14'b01_110100111110: DATA = 12'b100000000000;
            14'b01_110100111111: DATA = 12'b100000000000;
            14'b01_110101000000: DATA = 12'b100000000000;
            14'b01_110101000001: DATA = 12'b100000000000;
            14'b01_110101000010: DATA = 12'b100000000000;
            14'b01_110101000011: DATA = 12'b100000000000;
            14'b01_110101000100: DATA = 12'b100000000000;
            14'b01_110101000101: DATA = 12'b100000000000;
            14'b01_110101000110: DATA = 12'b100000000000;
            14'b01_110101000111: DATA = 12'b100000000000;
            14'b01_110101001000: DATA = 12'b100000000000;
            14'b01_110101001001: DATA = 12'b100000000000;
            14'b01_110101001010: DATA = 12'b100000000000;
            14'b01_110101001011: DATA = 12'b100000000000;
            14'b01_110101001100: DATA = 12'b100000000000;
            14'b01_110101001101: DATA = 12'b100000000000;
            14'b01_110101001110: DATA = 12'b100000000000;
            14'b01_110101001111: DATA = 12'b100000000000;
            14'b01_110101010000: DATA = 12'b100000000000;
            14'b01_110101010001: DATA = 12'b100000000000;
            14'b01_110101010010: DATA = 12'b100000000000;
            14'b01_110101010011: DATA = 12'b100000000000;
            14'b01_110101010100: DATA = 12'b100000000000;
            14'b01_110101010101: DATA = 12'b100000000000;
            14'b01_110101010110: DATA = 12'b100000000000;
            14'b01_110101010111: DATA = 12'b100000000000;
            14'b01_110101011000: DATA = 12'b100000000000;
            14'b01_110101011001: DATA = 12'b100000000000;
            14'b01_110101011010: DATA = 12'b100000000000;
            14'b01_110101011011: DATA = 12'b100000000000;
            14'b01_110101011100: DATA = 12'b100000000000;
            14'b01_110101011101: DATA = 12'b100000000000;
            14'b01_110101011110: DATA = 12'b100000000000;
            14'b01_110101011111: DATA = 12'b100000000000;
            14'b01_110101100000: DATA = 12'b100000000000;
            14'b01_110101100001: DATA = 12'b100000000000;
            14'b01_110101100010: DATA = 12'b100000000000;
            14'b01_110101100011: DATA = 12'b100000000000;
            14'b01_110101100100: DATA = 12'b100000000000;
            14'b01_110101100101: DATA = 12'b100000000000;
            14'b01_110101100110: DATA = 12'b100000000000;
            14'b01_110101100111: DATA = 12'b100000000000;
            14'b01_110101101000: DATA = 12'b100000000000;
            14'b01_110101101001: DATA = 12'b100000000000;
            14'b01_110101101010: DATA = 12'b100000000000;
            14'b01_110101101011: DATA = 12'b100000000000;
            14'b01_110101101100: DATA = 12'b100000000000;
            14'b01_110101101101: DATA = 12'b100000000000;
            14'b01_110101101110: DATA = 12'b100000000000;
            14'b01_110101101111: DATA = 12'b100000000000;
            14'b01_110101110000: DATA = 12'b100000000000;
            14'b01_110101110001: DATA = 12'b100000000000;
            14'b01_110101110010: DATA = 12'b100000000000;
            14'b01_110101110011: DATA = 12'b100000000000;
            14'b01_110101110100: DATA = 12'b100000000000;
            14'b01_110101110101: DATA = 12'b100000000000;
            14'b01_110101110110: DATA = 12'b100000000000;
            14'b01_110101110111: DATA = 12'b100000000000;
            14'b01_110101111000: DATA = 12'b100000000000;
            14'b01_110101111001: DATA = 12'b100000000000;
            14'b01_110101111010: DATA = 12'b100000000000;
            14'b01_110101111011: DATA = 12'b100000000000;
            14'b01_110101111100: DATA = 12'b100000000000;
            14'b01_110101111101: DATA = 12'b100000000000;
            14'b01_110101111110: DATA = 12'b100000000000;
            14'b01_110101111111: DATA = 12'b100000000000;
            14'b01_110110000000: DATA = 12'b100000000000;
            14'b01_110110000001: DATA = 12'b100000000000;
            14'b01_110110000010: DATA = 12'b100000000000;
            14'b01_110110000011: DATA = 12'b100000000000;
            14'b01_110110000100: DATA = 12'b100000000000;
            14'b01_110110000101: DATA = 12'b100000000000;
            14'b01_110110000110: DATA = 12'b100000000000;
            14'b01_110110000111: DATA = 12'b100000000000;
            14'b01_110110001000: DATA = 12'b100000000000;
            14'b01_110110001001: DATA = 12'b100000000000;
            14'b01_110110001010: DATA = 12'b100000000000;
            14'b01_110110001011: DATA = 12'b100000000000;
            14'b01_110110001100: DATA = 12'b100000000000;
            14'b01_110110001101: DATA = 12'b100000000000;
            14'b01_110110001110: DATA = 12'b100000000000;
            14'b01_110110001111: DATA = 12'b100000000000;
            14'b01_110110010000: DATA = 12'b100000000000;
            14'b01_110110010001: DATA = 12'b100000000000;
            14'b01_110110010010: DATA = 12'b100000000000;
            14'b01_110110010011: DATA = 12'b100000000000;
            14'b01_110110010100: DATA = 12'b100000000000;
            14'b01_110110010101: DATA = 12'b100000000000;
            14'b01_110110010110: DATA = 12'b100000000000;
            14'b01_110110010111: DATA = 12'b100000000000;
            14'b01_110110011000: DATA = 12'b100000000000;
            14'b01_110110011001: DATA = 12'b100000000000;
            14'b01_110110011010: DATA = 12'b100000000000;
            14'b01_110110011011: DATA = 12'b100000000000;
            14'b01_110110011100: DATA = 12'b100000000000;
            14'b01_110110011101: DATA = 12'b100000000000;
            14'b01_110110011110: DATA = 12'b100000000000;
            14'b01_110110011111: DATA = 12'b100000000000;
            14'b01_110110100000: DATA = 12'b100000000000;
            14'b01_110110100001: DATA = 12'b100000000000;
            14'b01_110110100010: DATA = 12'b100000000000;
            14'b01_110110100011: DATA = 12'b100000000000;
            14'b01_110110100100: DATA = 12'b100000000000;
            14'b01_110110100101: DATA = 12'b100000000000;
            14'b01_110110100110: DATA = 12'b100000000000;
            14'b01_110110100111: DATA = 12'b100000000000;
            14'b01_110110101000: DATA = 12'b100000000000;
            14'b01_110110101001: DATA = 12'b100000000000;
            14'b01_110110101010: DATA = 12'b100000000000;
            14'b01_110110101011: DATA = 12'b100000000000;
            14'b01_110110101100: DATA = 12'b100000000000;
            14'b01_110110101101: DATA = 12'b100000000000;
            14'b01_110110101110: DATA = 12'b100000000000;
            14'b01_110110101111: DATA = 12'b100000000000;
            14'b01_110110110000: DATA = 12'b100000000000;
            14'b01_110110110001: DATA = 12'b100000000000;
            14'b01_110110110010: DATA = 12'b100000000000;
            14'b01_110110110011: DATA = 12'b100000000000;
            14'b01_110110110100: DATA = 12'b100000000000;
            14'b01_110110110101: DATA = 12'b100000000000;
            14'b01_110110110110: DATA = 12'b100000000000;
            14'b01_110110110111: DATA = 12'b100000000000;
            14'b01_110110111000: DATA = 12'b100000000000;
            14'b01_110110111001: DATA = 12'b100000000000;
            14'b01_110110111010: DATA = 12'b100000000000;
            14'b01_110110111011: DATA = 12'b100000000000;
            14'b01_110110111100: DATA = 12'b100000000000;
            14'b01_110110111101: DATA = 12'b100000000000;
            14'b01_110110111110: DATA = 12'b100000000000;
            14'b01_110110111111: DATA = 12'b100000000000;
            14'b01_110111000000: DATA = 12'b100000000000;
            14'b01_110111000001: DATA = 12'b100000000000;
            14'b01_110111000010: DATA = 12'b100000000000;
            14'b01_110111000011: DATA = 12'b100000000000;
            14'b01_110111000100: DATA = 12'b100000000000;
            14'b01_110111000101: DATA = 12'b100000000000;
            14'b01_110111000110: DATA = 12'b100000000000;
            14'b01_110111000111: DATA = 12'b100000000000;
            14'b01_110111001000: DATA = 12'b100000000000;
            14'b01_110111001001: DATA = 12'b100000000000;
            14'b01_110111001010: DATA = 12'b100000000000;
            14'b01_110111001011: DATA = 12'b100000000000;
            14'b01_110111001100: DATA = 12'b100000000000;
            14'b01_110111001101: DATA = 12'b100000000000;
            14'b01_110111001110: DATA = 12'b100000000000;
            14'b01_110111001111: DATA = 12'b100000000000;
            14'b01_110111010000: DATA = 12'b100000000000;
            14'b01_110111010001: DATA = 12'b100000000000;
            14'b01_110111010010: DATA = 12'b100000000000;
            14'b01_110111010011: DATA = 12'b100000000000;
            14'b01_110111010100: DATA = 12'b100000000000;
            14'b01_110111010101: DATA = 12'b100000000000;
            14'b01_110111010110: DATA = 12'b100000000000;
            14'b01_110111010111: DATA = 12'b100000000000;
            14'b01_110111011000: DATA = 12'b100000000000;
            14'b01_110111011001: DATA = 12'b100000000000;
            14'b01_110111011010: DATA = 12'b100000000000;
            14'b01_110111011011: DATA = 12'b100000000000;
            14'b01_110111011100: DATA = 12'b100000000000;
            14'b01_110111011101: DATA = 12'b100000000000;
            14'b01_110111011110: DATA = 12'b100000000000;
            14'b01_110111011111: DATA = 12'b100000000000;
            14'b01_110111100000: DATA = 12'b100000000000;
            14'b01_110111100001: DATA = 12'b100000000000;
            14'b01_110111100010: DATA = 12'b100000000000;
            14'b01_110111100011: DATA = 12'b100000000000;
            14'b01_110111100100: DATA = 12'b100000000000;
            14'b01_110111100101: DATA = 12'b100000000000;
            14'b01_110111100110: DATA = 12'b100000000000;
            14'b01_110111100111: DATA = 12'b100000000000;
            14'b01_110111101000: DATA = 12'b100000000000;
            14'b01_110111101001: DATA = 12'b100000000000;
            14'b01_110111101010: DATA = 12'b100000000000;
            14'b01_110111101011: DATA = 12'b100000000000;
            14'b01_110111101100: DATA = 12'b100000000000;
            14'b01_110111101101: DATA = 12'b100000000000;
            14'b01_110111101110: DATA = 12'b100000000000;
            14'b01_110111101111: DATA = 12'b100000000000;
            14'b01_110111110000: DATA = 12'b100000000000;
            14'b01_110111110001: DATA = 12'b100000000000;
            14'b01_110111110010: DATA = 12'b100000000000;
            14'b01_110111110011: DATA = 12'b100000000000;
            14'b01_110111110100: DATA = 12'b100000000000;
            14'b01_110111110101: DATA = 12'b100000000000;
            14'b01_110111110110: DATA = 12'b100000000000;
            14'b01_110111110111: DATA = 12'b100000000000;
            14'b01_110111111000: DATA = 12'b100000000000;
            14'b01_110111111001: DATA = 12'b100000000000;
            14'b01_110111111010: DATA = 12'b100000000000;
            14'b01_110111111011: DATA = 12'b100000000000;
            14'b01_110111111100: DATA = 12'b100000000000;
            14'b01_110111111101: DATA = 12'b100000000000;
            14'b01_110111111110: DATA = 12'b100000000000;
            14'b01_110111111111: DATA = 12'b100000000000;
            14'b01_111000000000: DATA = 12'b100000000000;
            14'b01_111000000001: DATA = 12'b100000000000;
            14'b01_111000000010: DATA = 12'b100000000000;
            14'b01_111000000011: DATA = 12'b100000000000;
            14'b01_111000000100: DATA = 12'b100000000000;
            14'b01_111000000101: DATA = 12'b100000000000;
            14'b01_111000000110: DATA = 12'b100000000000;
            14'b01_111000000111: DATA = 12'b100000000000;
            14'b01_111000001000: DATA = 12'b100000000000;
            14'b01_111000001001: DATA = 12'b100000000000;
            14'b01_111000001010: DATA = 12'b100000000000;
            14'b01_111000001011: DATA = 12'b100000000000;
            14'b01_111000001100: DATA = 12'b100000000000;
            14'b01_111000001101: DATA = 12'b100000000000;
            14'b01_111000001110: DATA = 12'b100000000000;
            14'b01_111000001111: DATA = 12'b100000000000;
            14'b01_111000010000: DATA = 12'b100000000000;
            14'b01_111000010001: DATA = 12'b100000000000;
            14'b01_111000010010: DATA = 12'b100000000000;
            14'b01_111000010011: DATA = 12'b100000000000;
            14'b01_111000010100: DATA = 12'b100000000000;
            14'b01_111000010101: DATA = 12'b100000000000;
            14'b01_111000010110: DATA = 12'b100000000000;
            14'b01_111000010111: DATA = 12'b100000000000;
            14'b01_111000011000: DATA = 12'b100000000000;
            14'b01_111000011001: DATA = 12'b100000000000;
            14'b01_111000011010: DATA = 12'b100000000000;
            14'b01_111000011011: DATA = 12'b100000000000;
            14'b01_111000011100: DATA = 12'b100000000000;
            14'b01_111000011101: DATA = 12'b100000000000;
            14'b01_111000011110: DATA = 12'b100000000000;
            14'b01_111000011111: DATA = 12'b100000000000;
            14'b01_111000100000: DATA = 12'b100000000000;
            14'b01_111000100001: DATA = 12'b100000000000;
            14'b01_111000100010: DATA = 12'b100000000000;
            14'b01_111000100011: DATA = 12'b100000000000;
            14'b01_111000100100: DATA = 12'b100000000000;
            14'b01_111000100101: DATA = 12'b100000000000;
            14'b01_111000100110: DATA = 12'b100000000000;
            14'b01_111000100111: DATA = 12'b100000000000;
            14'b01_111000101000: DATA = 12'b100000000000;
            14'b01_111000101001: DATA = 12'b100000000000;
            14'b01_111000101010: DATA = 12'b100000000000;
            14'b01_111000101011: DATA = 12'b100000000000;
            14'b01_111000101100: DATA = 12'b100000000000;
            14'b01_111000101101: DATA = 12'b100000000000;
            14'b01_111000101110: DATA = 12'b100000000000;
            14'b01_111000101111: DATA = 12'b100000000000;
            14'b01_111000110000: DATA = 12'b100000000000;
            14'b01_111000110001: DATA = 12'b100000000000;
            14'b01_111000110010: DATA = 12'b100000000000;
            14'b01_111000110011: DATA = 12'b100000000000;
            14'b01_111000110100: DATA = 12'b100000000000;
            14'b01_111000110101: DATA = 12'b100000000000;
            14'b01_111000110110: DATA = 12'b100000000000;
            14'b01_111000110111: DATA = 12'b100000000000;
            14'b01_111000111000: DATA = 12'b100000000000;
            14'b01_111000111001: DATA = 12'b100000000000;
            14'b01_111000111010: DATA = 12'b100000000000;
            14'b01_111000111011: DATA = 12'b100000000000;
            14'b01_111000111100: DATA = 12'b100000000000;
            14'b01_111000111101: DATA = 12'b100000000000;
            14'b01_111000111110: DATA = 12'b100000000000;
            14'b01_111000111111: DATA = 12'b100000000000;
            14'b01_111001000000: DATA = 12'b100000000000;
            14'b01_111001000001: DATA = 12'b100000000000;
            14'b01_111001000010: DATA = 12'b100000000000;
            14'b01_111001000011: DATA = 12'b100000000000;
            14'b01_111001000100: DATA = 12'b100000000000;
            14'b01_111001000101: DATA = 12'b100000000000;
            14'b01_111001000110: DATA = 12'b100000000000;
            14'b01_111001000111: DATA = 12'b100000000000;
            14'b01_111001001000: DATA = 12'b100000000000;
            14'b01_111001001001: DATA = 12'b100000000000;
            14'b01_111001001010: DATA = 12'b100000000000;
            14'b01_111001001011: DATA = 12'b100000000000;
            14'b01_111001001100: DATA = 12'b100000000000;
            14'b01_111001001101: DATA = 12'b100000000000;
            14'b01_111001001110: DATA = 12'b100000000000;
            14'b01_111001001111: DATA = 12'b100000000000;
            14'b01_111001010000: DATA = 12'b100000000000;
            14'b01_111001010001: DATA = 12'b100000000000;
            14'b01_111001010010: DATA = 12'b100000000000;
            14'b01_111001010011: DATA = 12'b100000000000;
            14'b01_111001010100: DATA = 12'b100000000000;
            14'b01_111001010101: DATA = 12'b100000000000;
            14'b01_111001010110: DATA = 12'b100000000000;
            14'b01_111001010111: DATA = 12'b100000000000;
            14'b01_111001011000: DATA = 12'b100000000000;
            14'b01_111001011001: DATA = 12'b100000000000;
            14'b01_111001011010: DATA = 12'b100000000000;
            14'b01_111001011011: DATA = 12'b100000000000;
            14'b01_111001011100: DATA = 12'b100000000000;
            14'b01_111001011101: DATA = 12'b100000000000;
            14'b01_111001011110: DATA = 12'b100000000000;
            14'b01_111001011111: DATA = 12'b100000000000;
            14'b01_111001100000: DATA = 12'b100000000000;
            14'b01_111001100001: DATA = 12'b100000000000;
            14'b01_111001100010: DATA = 12'b100000000000;
            14'b01_111001100011: DATA = 12'b100000000000;
            14'b01_111001100100: DATA = 12'b100000000000;
            14'b01_111001100101: DATA = 12'b100000000000;
            14'b01_111001100110: DATA = 12'b100000000000;
            14'b01_111001100111: DATA = 12'b100000000000;
            14'b01_111001101000: DATA = 12'b100000000000;
            14'b01_111001101001: DATA = 12'b100000000000;
            14'b01_111001101010: DATA = 12'b100000000000;
            14'b01_111001101011: DATA = 12'b100000000000;
            14'b01_111001101100: DATA = 12'b100000000000;
            14'b01_111001101101: DATA = 12'b100000000000;
            14'b01_111001101110: DATA = 12'b100000000000;
            14'b01_111001101111: DATA = 12'b100000000000;
            14'b01_111001110000: DATA = 12'b100000000000;
            14'b01_111001110001: DATA = 12'b100000000000;
            14'b01_111001110010: DATA = 12'b100000000000;
            14'b01_111001110011: DATA = 12'b100000000000;
            14'b01_111001110100: DATA = 12'b100000000000;
            14'b01_111001110101: DATA = 12'b100000000000;
            14'b01_111001110110: DATA = 12'b100000000000;
            14'b01_111001110111: DATA = 12'b100000000000;
            14'b01_111001111000: DATA = 12'b100000000000;
            14'b01_111001111001: DATA = 12'b100000000000;
            14'b01_111001111010: DATA = 12'b100000000000;
            14'b01_111001111011: DATA = 12'b100000000000;
            14'b01_111001111100: DATA = 12'b100000000000;
            14'b01_111001111101: DATA = 12'b100000000000;
            14'b01_111001111110: DATA = 12'b100000000000;
            14'b01_111001111111: DATA = 12'b100000000000;
            14'b01_111010000000: DATA = 12'b100000000000;
            14'b01_111010000001: DATA = 12'b100000000000;
            14'b01_111010000010: DATA = 12'b100000000000;
            14'b01_111010000011: DATA = 12'b100000000000;
            14'b01_111010000100: DATA = 12'b100000000000;
            14'b01_111010000101: DATA = 12'b100000000000;
            14'b01_111010000110: DATA = 12'b100000000000;
            14'b01_111010000111: DATA = 12'b100000000000;
            14'b01_111010001000: DATA = 12'b100000000000;
            14'b01_111010001001: DATA = 12'b100000000000;
            14'b01_111010001010: DATA = 12'b100000000000;
            14'b01_111010001011: DATA = 12'b100000000000;
            14'b01_111010001100: DATA = 12'b100000000000;
            14'b01_111010001101: DATA = 12'b100000000000;
            14'b01_111010001110: DATA = 12'b100000000000;
            14'b01_111010001111: DATA = 12'b100000000000;
            14'b01_111010010000: DATA = 12'b100000000000;
            14'b01_111010010001: DATA = 12'b100000000000;
            14'b01_111010010010: DATA = 12'b100000000000;
            14'b01_111010010011: DATA = 12'b100000000000;
            14'b01_111010010100: DATA = 12'b100000000000;
            14'b01_111010010101: DATA = 12'b100000000000;
            14'b01_111010010110: DATA = 12'b100000000000;
            14'b01_111010010111: DATA = 12'b100000000000;
            14'b01_111010011000: DATA = 12'b100000000000;
            14'b01_111010011001: DATA = 12'b100000000000;
            14'b01_111010011010: DATA = 12'b100000000000;
            14'b01_111010011011: DATA = 12'b100000000000;
            14'b01_111010011100: DATA = 12'b100000000000;
            14'b01_111010011101: DATA = 12'b100000000000;
            14'b01_111010011110: DATA = 12'b100000000000;
            14'b01_111010011111: DATA = 12'b100000000000;
            14'b01_111010100000: DATA = 12'b100000000000;
            14'b01_111010100001: DATA = 12'b100000000000;
            14'b01_111010100010: DATA = 12'b100000000000;
            14'b01_111010100011: DATA = 12'b100000000000;
            14'b01_111010100100: DATA = 12'b100000000000;
            14'b01_111010100101: DATA = 12'b100000000000;
            14'b01_111010100110: DATA = 12'b100000000000;
            14'b01_111010100111: DATA = 12'b100000000000;
            14'b01_111010101000: DATA = 12'b100000000000;
            14'b01_111010101001: DATA = 12'b100000000000;
            14'b01_111010101010: DATA = 12'b100000000000;
            14'b01_111010101011: DATA = 12'b100000000000;
            14'b01_111010101100: DATA = 12'b100000000000;
            14'b01_111010101101: DATA = 12'b100000000000;
            14'b01_111010101110: DATA = 12'b100000000000;
            14'b01_111010101111: DATA = 12'b100000000000;
            14'b01_111010110000: DATA = 12'b100000000000;
            14'b01_111010110001: DATA = 12'b100000000000;
            14'b01_111010110010: DATA = 12'b100000000000;
            14'b01_111010110011: DATA = 12'b100000000000;
            14'b01_111010110100: DATA = 12'b100000000000;
            14'b01_111010110101: DATA = 12'b100000000000;
            14'b01_111010110110: DATA = 12'b100000000000;
            14'b01_111010110111: DATA = 12'b100000000000;
            14'b01_111010111000: DATA = 12'b100000000000;
            14'b01_111010111001: DATA = 12'b100000000000;
            14'b01_111010111010: DATA = 12'b100000000000;
            14'b01_111010111011: DATA = 12'b100000000000;
            14'b01_111010111100: DATA = 12'b100000000000;
            14'b01_111010111101: DATA = 12'b100000000000;
            14'b01_111010111110: DATA = 12'b100000000000;
            14'b01_111010111111: DATA = 12'b100000000000;
            14'b01_111011000000: DATA = 12'b100000000000;
            14'b01_111011000001: DATA = 12'b100000000000;
            14'b01_111011000010: DATA = 12'b100000000000;
            14'b01_111011000011: DATA = 12'b100000000000;
            14'b01_111011000100: DATA = 12'b100000000000;
            14'b01_111011000101: DATA = 12'b100000000000;
            14'b01_111011000110: DATA = 12'b100000000000;
            14'b01_111011000111: DATA = 12'b100000000000;
            14'b01_111011001000: DATA = 12'b100000000000;
            14'b01_111011001001: DATA = 12'b100000000000;
            14'b01_111011001010: DATA = 12'b100000000000;
            14'b01_111011001011: DATA = 12'b100000000000;
            14'b01_111011001100: DATA = 12'b100000000000;
            14'b01_111011001101: DATA = 12'b100000000000;
            14'b01_111011001110: DATA = 12'b100000000000;
            14'b01_111011001111: DATA = 12'b100000000000;
            14'b01_111011010000: DATA = 12'b100000000000;
            14'b01_111011010001: DATA = 12'b100000000000;
            14'b01_111011010010: DATA = 12'b100000000000;
            14'b01_111011010011: DATA = 12'b100000000000;
            14'b01_111011010100: DATA = 12'b100000000000;
            14'b01_111011010101: DATA = 12'b100000000000;
            14'b01_111011010110: DATA = 12'b100000000000;
            14'b01_111011010111: DATA = 12'b100000000000;
            14'b01_111011011000: DATA = 12'b100000000000;
            14'b01_111011011001: DATA = 12'b100000000000;
            14'b01_111011011010: DATA = 12'b100000000000;
            14'b01_111011011011: DATA = 12'b100000000000;
            14'b01_111011011100: DATA = 12'b100000000000;
            14'b01_111011011101: DATA = 12'b100000000000;
            14'b01_111011011110: DATA = 12'b100000000000;
            14'b01_111011011111: DATA = 12'b100000000000;
            14'b01_111011100000: DATA = 12'b100000000000;
            14'b01_111011100001: DATA = 12'b100000000000;
            14'b01_111011100010: DATA = 12'b100000000000;
            14'b01_111011100011: DATA = 12'b100000000000;
            14'b01_111011100100: DATA = 12'b100000000000;
            14'b01_111011100101: DATA = 12'b100000000000;
            14'b01_111011100110: DATA = 12'b100000000000;
            14'b01_111011100111: DATA = 12'b100000000000;
            14'b01_111011101000: DATA = 12'b100000000000;
            14'b01_111011101001: DATA = 12'b100000000000;
            14'b01_111011101010: DATA = 12'b100000000000;
            14'b01_111011101011: DATA = 12'b100000000000;
            14'b01_111011101100: DATA = 12'b100000000000;
            14'b01_111011101101: DATA = 12'b100000000000;
            14'b01_111011101110: DATA = 12'b100000000000;
            14'b01_111011101111: DATA = 12'b100000000000;
            14'b01_111011110000: DATA = 12'b100000000000;
            14'b01_111011110001: DATA = 12'b100000000000;
            14'b01_111011110010: DATA = 12'b100000000000;
            14'b01_111011110011: DATA = 12'b100000000000;
            14'b01_111011110100: DATA = 12'b100000000000;
            14'b01_111011110101: DATA = 12'b100000000000;
            14'b01_111011110110: DATA = 12'b100000000000;
            14'b01_111011110111: DATA = 12'b100000000000;
            14'b01_111011111000: DATA = 12'b100000000000;
            14'b01_111011111001: DATA = 12'b100000000000;
            14'b01_111011111010: DATA = 12'b100000000000;
            14'b01_111011111011: DATA = 12'b100000000000;
            14'b01_111011111100: DATA = 12'b100000000000;
            14'b01_111011111101: DATA = 12'b100000000000;
            14'b01_111011111110: DATA = 12'b100000000000;
            14'b01_111011111111: DATA = 12'b100000000000;
            14'b01_111100000000: DATA = 12'b100000000000;
            14'b01_111100000001: DATA = 12'b100000000000;
            14'b01_111100000010: DATA = 12'b100000000000;
            14'b01_111100000011: DATA = 12'b100000000000;
            14'b01_111100000100: DATA = 12'b100000000000;
            14'b01_111100000101: DATA = 12'b100000000000;
            14'b01_111100000110: DATA = 12'b100000000000;
            14'b01_111100000111: DATA = 12'b100000000000;
            14'b01_111100001000: DATA = 12'b100000000000;
            14'b01_111100001001: DATA = 12'b100000000000;
            14'b01_111100001010: DATA = 12'b100000000000;
            14'b01_111100001011: DATA = 12'b100000000000;
            14'b01_111100001100: DATA = 12'b100000000000;
            14'b01_111100001101: DATA = 12'b100000000000;
            14'b01_111100001110: DATA = 12'b100000000000;
            14'b01_111100001111: DATA = 12'b100000000000;
            14'b01_111100010000: DATA = 12'b100000000000;
            14'b01_111100010001: DATA = 12'b100000000000;
            14'b01_111100010010: DATA = 12'b100000000000;
            14'b01_111100010011: DATA = 12'b100000000000;
            14'b01_111100010100: DATA = 12'b100000000000;
            14'b01_111100010101: DATA = 12'b100000000000;
            14'b01_111100010110: DATA = 12'b100000000000;
            14'b01_111100010111: DATA = 12'b100000000000;
            14'b01_111100011000: DATA = 12'b100000000000;
            14'b01_111100011001: DATA = 12'b100000000000;
            14'b01_111100011010: DATA = 12'b100000000000;
            14'b01_111100011011: DATA = 12'b100000000000;
            14'b01_111100011100: DATA = 12'b100000000000;
            14'b01_111100011101: DATA = 12'b100000000000;
            14'b01_111100011110: DATA = 12'b100000000000;
            14'b01_111100011111: DATA = 12'b100000000000;
            14'b01_111100100000: DATA = 12'b100000000000;
            14'b01_111100100001: DATA = 12'b100000000000;
            14'b01_111100100010: DATA = 12'b100000000000;
            14'b01_111100100011: DATA = 12'b100000000000;
            14'b01_111100100100: DATA = 12'b100000000000;
            14'b01_111100100101: DATA = 12'b100000000000;
            14'b01_111100100110: DATA = 12'b100000000000;
            14'b01_111100100111: DATA = 12'b100000000000;
            14'b01_111100101000: DATA = 12'b100000000000;
            14'b01_111100101001: DATA = 12'b100000000000;
            14'b01_111100101010: DATA = 12'b100000000000;
            14'b01_111100101011: DATA = 12'b100000000000;
            14'b01_111100101100: DATA = 12'b100000000000;
            14'b01_111100101101: DATA = 12'b100000000000;
            14'b01_111100101110: DATA = 12'b100000000000;
            14'b01_111100101111: DATA = 12'b100000000000;
            14'b01_111100110000: DATA = 12'b100000000000;
            14'b01_111100110001: DATA = 12'b100000000000;
            14'b01_111100110010: DATA = 12'b100000000000;
            14'b01_111100110011: DATA = 12'b100000000000;
            14'b01_111100110100: DATA = 12'b100000000000;
            14'b01_111100110101: DATA = 12'b100000000000;
            14'b01_111100110110: DATA = 12'b100000000000;
            14'b01_111100110111: DATA = 12'b100000000000;
            14'b01_111100111000: DATA = 12'b100000000000;
            14'b01_111100111001: DATA = 12'b100000000000;
            14'b01_111100111010: DATA = 12'b100000000000;
            14'b01_111100111011: DATA = 12'b100000000000;
            14'b01_111100111100: DATA = 12'b100000000000;
            14'b01_111100111101: DATA = 12'b100000000000;
            14'b01_111100111110: DATA = 12'b100000000000;
            14'b01_111100111111: DATA = 12'b100000000000;
            14'b01_111101000000: DATA = 12'b100000000000;
            14'b01_111101000001: DATA = 12'b100000000000;
            14'b01_111101000010: DATA = 12'b100000000000;
            14'b01_111101000011: DATA = 12'b100000000000;
            14'b01_111101000100: DATA = 12'b100000000000;
            14'b01_111101000101: DATA = 12'b100000000000;
            14'b01_111101000110: DATA = 12'b100000000000;
            14'b01_111101000111: DATA = 12'b100000000000;
            14'b01_111101001000: DATA = 12'b100000000000;
            14'b01_111101001001: DATA = 12'b100000000000;
            14'b01_111101001010: DATA = 12'b100000000000;
            14'b01_111101001011: DATA = 12'b100000000000;
            14'b01_111101001100: DATA = 12'b100000000000;
            14'b01_111101001101: DATA = 12'b100000000000;
            14'b01_111101001110: DATA = 12'b100000000000;
            14'b01_111101001111: DATA = 12'b100000000000;
            14'b01_111101010000: DATA = 12'b100000000000;
            14'b01_111101010001: DATA = 12'b100000000000;
            14'b01_111101010010: DATA = 12'b100000000000;
            14'b01_111101010011: DATA = 12'b100000000000;
            14'b01_111101010100: DATA = 12'b100000000000;
            14'b01_111101010101: DATA = 12'b100000000000;
            14'b01_111101010110: DATA = 12'b100000000000;
            14'b01_111101010111: DATA = 12'b100000000000;
            14'b01_111101011000: DATA = 12'b100000000000;
            14'b01_111101011001: DATA = 12'b100000000000;
            14'b01_111101011010: DATA = 12'b100000000000;
            14'b01_111101011011: DATA = 12'b100000000000;
            14'b01_111101011100: DATA = 12'b100000000000;
            14'b01_111101011101: DATA = 12'b100000000000;
            14'b01_111101011110: DATA = 12'b100000000000;
            14'b01_111101011111: DATA = 12'b100000000000;
            14'b01_111101100000: DATA = 12'b100000000000;
            14'b01_111101100001: DATA = 12'b100000000000;
            14'b01_111101100010: DATA = 12'b100000000000;
            14'b01_111101100011: DATA = 12'b100000000000;
            14'b01_111101100100: DATA = 12'b100000000000;
            14'b01_111101100101: DATA = 12'b100000000000;
            14'b01_111101100110: DATA = 12'b100000000000;
            14'b01_111101100111: DATA = 12'b100000000000;
            14'b01_111101101000: DATA = 12'b100000000000;
            14'b01_111101101001: DATA = 12'b100000000000;
            14'b01_111101101010: DATA = 12'b100000000000;
            14'b01_111101101011: DATA = 12'b100000000000;
            14'b01_111101101100: DATA = 12'b100000000000;
            14'b01_111101101101: DATA = 12'b100000000000;
            14'b01_111101101110: DATA = 12'b100000000000;
            14'b01_111101101111: DATA = 12'b100000000000;
            14'b01_111101110000: DATA = 12'b100000000000;
            14'b01_111101110001: DATA = 12'b100000000000;
            14'b01_111101110010: DATA = 12'b100000000000;
            14'b01_111101110011: DATA = 12'b100000000000;
            14'b01_111101110100: DATA = 12'b100000000000;
            14'b01_111101110101: DATA = 12'b100000000000;
            14'b01_111101110110: DATA = 12'b100000000000;
            14'b01_111101110111: DATA = 12'b100000000000;
            14'b01_111101111000: DATA = 12'b100000000000;
            14'b01_111101111001: DATA = 12'b100000000000;
            14'b01_111101111010: DATA = 12'b100000000000;
            14'b01_111101111011: DATA = 12'b100000000000;
            14'b01_111101111100: DATA = 12'b100000000000;
            14'b01_111101111101: DATA = 12'b100000000000;
            14'b01_111101111110: DATA = 12'b100000000000;
            14'b01_111101111111: DATA = 12'b100000000000;
            14'b01_111110000000: DATA = 12'b100000000000;
            14'b01_111110000001: DATA = 12'b100000000000;
            14'b01_111110000010: DATA = 12'b100000000000;
            14'b01_111110000011: DATA = 12'b100000000000;
            14'b01_111110000100: DATA = 12'b100000000000;
            14'b01_111110000101: DATA = 12'b100000000000;
            14'b01_111110000110: DATA = 12'b100000000000;
            14'b01_111110000111: DATA = 12'b100000000000;
            14'b01_111110001000: DATA = 12'b100000000000;
            14'b01_111110001001: DATA = 12'b100000000000;
            14'b01_111110001010: DATA = 12'b100000000000;
            14'b01_111110001011: DATA = 12'b100000000000;
            14'b01_111110001100: DATA = 12'b100000000000;
            14'b01_111110001101: DATA = 12'b100000000000;
            14'b01_111110001110: DATA = 12'b100000000000;
            14'b01_111110001111: DATA = 12'b100000000000;
            14'b01_111110010000: DATA = 12'b100000000000;
            14'b01_111110010001: DATA = 12'b100000000000;
            14'b01_111110010010: DATA = 12'b100000000000;
            14'b01_111110010011: DATA = 12'b100000000000;
            14'b01_111110010100: DATA = 12'b100000000000;
            14'b01_111110010101: DATA = 12'b100000000000;
            14'b01_111110010110: DATA = 12'b100000000000;
            14'b01_111110010111: DATA = 12'b100000000000;
            14'b01_111110011000: DATA = 12'b100000000000;
            14'b01_111110011001: DATA = 12'b100000000000;
            14'b01_111110011010: DATA = 12'b100000000000;
            14'b01_111110011011: DATA = 12'b100000000000;
            14'b01_111110011100: DATA = 12'b100000000000;
            14'b01_111110011101: DATA = 12'b100000000000;
            14'b01_111110011110: DATA = 12'b100000000000;
            14'b01_111110011111: DATA = 12'b100000000000;
            14'b01_111110100000: DATA = 12'b100000000000;
            14'b01_111110100001: DATA = 12'b100000000000;
            14'b01_111110100010: DATA = 12'b100000000000;
            14'b01_111110100011: DATA = 12'b100000000000;
            14'b01_111110100100: DATA = 12'b100000000000;
            14'b01_111110100101: DATA = 12'b100000000000;
            14'b01_111110100110: DATA = 12'b100000000000;
            14'b01_111110100111: DATA = 12'b100000000000;
            14'b01_111110101000: DATA = 12'b100000000000;
            14'b01_111110101001: DATA = 12'b100000000000;
            14'b01_111110101010: DATA = 12'b100000000000;
            14'b01_111110101011: DATA = 12'b100000000000;
            14'b01_111110101100: DATA = 12'b100000000000;
            14'b01_111110101101: DATA = 12'b100000000000;
            14'b01_111110101110: DATA = 12'b100000000000;
            14'b01_111110101111: DATA = 12'b100000000000;
            14'b01_111110110000: DATA = 12'b100000000000;
            14'b01_111110110001: DATA = 12'b100000000000;
            14'b01_111110110010: DATA = 12'b100000000000;
            14'b01_111110110011: DATA = 12'b100000000000;
            14'b01_111110110100: DATA = 12'b100000000000;
            14'b01_111110110101: DATA = 12'b100000000000;
            14'b01_111110110110: DATA = 12'b100000000000;
            14'b01_111110110111: DATA = 12'b100000000000;
            14'b01_111110111000: DATA = 12'b100000000000;
            14'b01_111110111001: DATA = 12'b100000000000;
            14'b01_111110111010: DATA = 12'b100000000000;
            14'b01_111110111011: DATA = 12'b100000000000;
            14'b01_111110111100: DATA = 12'b100000000000;
            14'b01_111110111101: DATA = 12'b100000000000;
            14'b01_111110111110: DATA = 12'b100000000000;
            14'b01_111110111111: DATA = 12'b100000000000;
            14'b01_111111000000: DATA = 12'b100000000000;
            14'b01_111111000001: DATA = 12'b100000000000;
            14'b01_111111000010: DATA = 12'b100000000000;
            14'b01_111111000011: DATA = 12'b100000000000;
            14'b01_111111000100: DATA = 12'b100000000000;
            14'b01_111111000101: DATA = 12'b100000000000;
            14'b01_111111000110: DATA = 12'b100000000000;
            14'b01_111111000111: DATA = 12'b100000000000;
            14'b01_111111001000: DATA = 12'b100000000000;
            14'b01_111111001001: DATA = 12'b100000000000;
            14'b01_111111001010: DATA = 12'b100000000000;
            14'b01_111111001011: DATA = 12'b100000000000;
            14'b01_111111001100: DATA = 12'b100000000000;
            14'b01_111111001101: DATA = 12'b100000000000;
            14'b01_111111001110: DATA = 12'b100000000000;
            14'b01_111111001111: DATA = 12'b100000000000;
            14'b01_111111010000: DATA = 12'b100000000000;
            14'b01_111111010001: DATA = 12'b100000000000;
            14'b01_111111010010: DATA = 12'b100000000000;
            14'b01_111111010011: DATA = 12'b100000000000;
            14'b01_111111010100: DATA = 12'b100000000000;
            14'b01_111111010101: DATA = 12'b100000000000;
            14'b01_111111010110: DATA = 12'b100000000000;
            14'b01_111111010111: DATA = 12'b100000000000;
            14'b01_111111011000: DATA = 12'b100000000000;
            14'b01_111111011001: DATA = 12'b100000000000;
            14'b01_111111011010: DATA = 12'b100000000000;
            14'b01_111111011011: DATA = 12'b100000000000;
            14'b01_111111011100: DATA = 12'b100000000000;
            14'b01_111111011101: DATA = 12'b100000000000;
            14'b01_111111011110: DATA = 12'b100000000000;
            14'b01_111111011111: DATA = 12'b100000000000;
            14'b01_111111100000: DATA = 12'b100000000000;
            14'b01_111111100001: DATA = 12'b100000000000;
            14'b01_111111100010: DATA = 12'b100000000000;
            14'b01_111111100011: DATA = 12'b100000000000;
            14'b01_111111100100: DATA = 12'b100000000000;
            14'b01_111111100101: DATA = 12'b100000000000;
            14'b01_111111100110: DATA = 12'b100000000000;
            14'b01_111111100111: DATA = 12'b100000000000;
            14'b01_111111101000: DATA = 12'b100000000000;
            14'b01_111111101001: DATA = 12'b100000000000;
            14'b01_111111101010: DATA = 12'b100000000000;
            14'b01_111111101011: DATA = 12'b100000000000;
            14'b01_111111101100: DATA = 12'b100000000000;
            14'b01_111111101101: DATA = 12'b100000000000;
            14'b01_111111101110: DATA = 12'b100000000000;
            14'b01_111111101111: DATA = 12'b100000000000;
            14'b01_111111110000: DATA = 12'b100000000000;
            14'b01_111111110001: DATA = 12'b100000000000;
            14'b01_111111110010: DATA = 12'b100000000000;
            14'b01_111111110011: DATA = 12'b100000000000;
            14'b01_111111110100: DATA = 12'b100000000000;
            14'b01_111111110101: DATA = 12'b100000000000;
            14'b01_111111110110: DATA = 12'b100000000000;
            14'b01_111111110111: DATA = 12'b100000000000;
            14'b01_111111111000: DATA = 12'b100000000000;
            14'b01_111111111001: DATA = 12'b100000000000;
            14'b01_111111111010: DATA = 12'b100000000000;
            14'b01_111111111011: DATA = 12'b100000000000;
            14'b01_111111111100: DATA = 12'b100000000000;
            14'b01_111111111101: DATA = 12'b100000000000;
            14'b01_111111111110: DATA = 12'b100000000000;
            14'b01_111111111111: DATA = 12'b100000000000;
            14'b10_000000000000: DATA = 12'b100000000000;
            14'b10_000000000001: DATA = 12'b011111111100;
            14'b10_000000000010: DATA = 12'b011111111001;
            14'b10_000000000011: DATA = 12'b011111110110;
            14'b10_000000000100: DATA = 12'b011111110011;
            14'b10_000000000101: DATA = 12'b011111110000;
            14'b10_000000000110: DATA = 12'b011111101101;
            14'b10_000000000111: DATA = 12'b011111101010;
            14'b10_000000001000: DATA = 12'b011111100110;
            14'b10_000000001001: DATA = 12'b011111100011;
            14'b10_000000001010: DATA = 12'b011111100000;
            14'b10_000000001011: DATA = 12'b011111011101;
            14'b10_000000001100: DATA = 12'b011111011010;
            14'b10_000000001101: DATA = 12'b011111010111;
            14'b10_000000001110: DATA = 12'b011111010100;
            14'b10_000000001111: DATA = 12'b011111010000;
            14'b10_000000010000: DATA = 12'b011111001101;
            14'b10_000000010001: DATA = 12'b011111001010;
            14'b10_000000010010: DATA = 12'b011111000111;
            14'b10_000000010011: DATA = 12'b011111000100;
            14'b10_000000010100: DATA = 12'b011111000001;
            14'b10_000000010101: DATA = 12'b011110111110;
            14'b10_000000010110: DATA = 12'b011110111010;
            14'b10_000000010111: DATA = 12'b011110110111;
            14'b10_000000011000: DATA = 12'b011110110100;
            14'b10_000000011001: DATA = 12'b011110110001;
            14'b10_000000011010: DATA = 12'b011110101110;
            14'b10_000000011011: DATA = 12'b011110101011;
            14'b10_000000011100: DATA = 12'b011110101000;
            14'b10_000000011101: DATA = 12'b011110100100;
            14'b10_000000011110: DATA = 12'b011110100001;
            14'b10_000000011111: DATA = 12'b011110011110;
            14'b10_000000100000: DATA = 12'b011110011011;
            14'b10_000000100001: DATA = 12'b011110011000;
            14'b10_000000100010: DATA = 12'b011110010101;
            14'b10_000000100011: DATA = 12'b011110010010;
            14'b10_000000100100: DATA = 12'b011110001111;
            14'b10_000000100101: DATA = 12'b011110001011;
            14'b10_000000100110: DATA = 12'b011110001000;
            14'b10_000000100111: DATA = 12'b011110000101;
            14'b10_000000101000: DATA = 12'b011110000010;
            14'b10_000000101001: DATA = 12'b011101111111;
            14'b10_000000101010: DATA = 12'b011101111100;
            14'b10_000000101011: DATA = 12'b011101111001;
            14'b10_000000101100: DATA = 12'b011101110101;
            14'b10_000000101101: DATA = 12'b011101110010;
            14'b10_000000101110: DATA = 12'b011101101111;
            14'b10_000000101111: DATA = 12'b011101101100;
            14'b10_000000110000: DATA = 12'b011101101001;
            14'b10_000000110001: DATA = 12'b011101100110;
            14'b10_000000110010: DATA = 12'b011101100011;
            14'b10_000000110011: DATA = 12'b011101100000;
            14'b10_000000110100: DATA = 12'b011101011100;
            14'b10_000000110101: DATA = 12'b011101011001;
            14'b10_000000110110: DATA = 12'b011101010110;
            14'b10_000000110111: DATA = 12'b011101010011;
            14'b10_000000111000: DATA = 12'b011101010000;
            14'b10_000000111001: DATA = 12'b011101001101;
            14'b10_000000111010: DATA = 12'b011101001010;
            14'b10_000000111011: DATA = 12'b011101000110;
            14'b10_000000111100: DATA = 12'b011101000011;
            14'b10_000000111101: DATA = 12'b011101000000;
            14'b10_000000111110: DATA = 12'b011100111101;
            14'b10_000000111111: DATA = 12'b011100111010;
            14'b10_000001000000: DATA = 12'b011100110111;
            14'b10_000001000001: DATA = 12'b011100110100;
            14'b10_000001000010: DATA = 12'b011100110001;
            14'b10_000001000011: DATA = 12'b011100101101;
            14'b10_000001000100: DATA = 12'b011100101010;
            14'b10_000001000101: DATA = 12'b011100100111;
            14'b10_000001000110: DATA = 12'b011100100100;
            14'b10_000001000111: DATA = 12'b011100100001;
            14'b10_000001001000: DATA = 12'b011100011110;
            14'b10_000001001001: DATA = 12'b011100011011;
            14'b10_000001001010: DATA = 12'b011100011000;
            14'b10_000001001011: DATA = 12'b011100010101;
            14'b10_000001001100: DATA = 12'b011100010001;
            14'b10_000001001101: DATA = 12'b011100001110;
            14'b10_000001001110: DATA = 12'b011100001011;
            14'b10_000001001111: DATA = 12'b011100001000;
            14'b10_000001010000: DATA = 12'b011100000101;
            14'b10_000001010001: DATA = 12'b011100000010;
            14'b10_000001010010: DATA = 12'b011011111111;
            14'b10_000001010011: DATA = 12'b011011111100;
            14'b10_000001010100: DATA = 12'b011011111000;
            14'b10_000001010101: DATA = 12'b011011110101;
            14'b10_000001010110: DATA = 12'b011011110010;
            14'b10_000001010111: DATA = 12'b011011101111;
            14'b10_000001011000: DATA = 12'b011011101100;
            14'b10_000001011001: DATA = 12'b011011101001;
            14'b10_000001011010: DATA = 12'b011011100110;
            14'b10_000001011011: DATA = 12'b011011100011;
            14'b10_000001011100: DATA = 12'b011011100000;
            14'b10_000001011101: DATA = 12'b011011011100;
            14'b10_000001011110: DATA = 12'b011011011001;
            14'b10_000001011111: DATA = 12'b011011010110;
            14'b10_000001100000: DATA = 12'b011011010011;
            14'b10_000001100001: DATA = 12'b011011010000;
            14'b10_000001100010: DATA = 12'b011011001101;
            14'b10_000001100011: DATA = 12'b011011001010;
            14'b10_000001100100: DATA = 12'b011011000111;
            14'b10_000001100101: DATA = 12'b011011000100;
            14'b10_000001100110: DATA = 12'b011011000001;
            14'b10_000001100111: DATA = 12'b011010111101;
            14'b10_000001101000: DATA = 12'b011010111010;
            14'b10_000001101001: DATA = 12'b011010110111;
            14'b10_000001101010: DATA = 12'b011010110100;
            14'b10_000001101011: DATA = 12'b011010110001;
            14'b10_000001101100: DATA = 12'b011010101110;
            14'b10_000001101101: DATA = 12'b011010101011;
            14'b10_000001101110: DATA = 12'b011010101000;
            14'b10_000001101111: DATA = 12'b011010100101;
            14'b10_000001110000: DATA = 12'b011010100010;
            14'b10_000001110001: DATA = 12'b011010011110;
            14'b10_000001110010: DATA = 12'b011010011011;
            14'b10_000001110011: DATA = 12'b011010011000;
            14'b10_000001110100: DATA = 12'b011010010101;
            14'b10_000001110101: DATA = 12'b011010010010;
            14'b10_000001110110: DATA = 12'b011010001111;
            14'b10_000001110111: DATA = 12'b011010001100;
            14'b10_000001111000: DATA = 12'b011010001001;
            14'b10_000001111001: DATA = 12'b011010000110;
            14'b10_000001111010: DATA = 12'b011010000011;
            14'b10_000001111011: DATA = 12'b011010000000;
            14'b10_000001111100: DATA = 12'b011001111100;
            14'b10_000001111101: DATA = 12'b011001111001;
            14'b10_000001111110: DATA = 12'b011001110110;
            14'b10_000001111111: DATA = 12'b011001110011;
            14'b10_000010000000: DATA = 12'b011001110000;
            14'b10_000010000001: DATA = 12'b011001101101;
            14'b10_000010000010: DATA = 12'b011001101010;
            14'b10_000010000011: DATA = 12'b011001100111;
            14'b10_000010000100: DATA = 12'b011001100100;
            14'b10_000010000101: DATA = 12'b011001100001;
            14'b10_000010000110: DATA = 12'b011001011110;
            14'b10_000010000111: DATA = 12'b011001011011;
            14'b10_000010001000: DATA = 12'b011001011000;
            14'b10_000010001001: DATA = 12'b011001010100;
            14'b10_000010001010: DATA = 12'b011001010001;
            14'b10_000010001011: DATA = 12'b011001001110;
            14'b10_000010001100: DATA = 12'b011001001011;
            14'b10_000010001101: DATA = 12'b011001001000;
            14'b10_000010001110: DATA = 12'b011001000101;
            14'b10_000010001111: DATA = 12'b011001000010;
            14'b10_000010010000: DATA = 12'b011000111111;
            14'b10_000010010001: DATA = 12'b011000111100;
            14'b10_000010010010: DATA = 12'b011000111001;
            14'b10_000010010011: DATA = 12'b011000110110;
            14'b10_000010010100: DATA = 12'b011000110011;
            14'b10_000010010101: DATA = 12'b011000110000;
            14'b10_000010010110: DATA = 12'b011000101101;
            14'b10_000010010111: DATA = 12'b011000101010;
            14'b10_000010011000: DATA = 12'b011000100111;
            14'b10_000010011001: DATA = 12'b011000100011;
            14'b10_000010011010: DATA = 12'b011000100000;
            14'b10_000010011011: DATA = 12'b011000011101;
            14'b10_000010011100: DATA = 12'b011000011010;
            14'b10_000010011101: DATA = 12'b011000010111;
            14'b10_000010011110: DATA = 12'b011000010100;
            14'b10_000010011111: DATA = 12'b011000010001;
            14'b10_000010100000: DATA = 12'b011000001110;
            14'b10_000010100001: DATA = 12'b011000001011;
            14'b10_000010100010: DATA = 12'b011000001000;
            14'b10_000010100011: DATA = 12'b011000000101;
            14'b10_000010100100: DATA = 12'b011000000010;
            14'b10_000010100101: DATA = 12'b010111111111;
            14'b10_000010100110: DATA = 12'b010111111100;
            14'b10_000010100111: DATA = 12'b010111111001;
            14'b10_000010101000: DATA = 12'b010111110110;
            14'b10_000010101001: DATA = 12'b010111110011;
            14'b10_000010101010: DATA = 12'b010111110000;
            14'b10_000010101011: DATA = 12'b010111101101;
            14'b10_000010101100: DATA = 12'b010111101010;
            14'b10_000010101101: DATA = 12'b010111100111;
            14'b10_000010101110: DATA = 12'b010111100100;
            14'b10_000010101111: DATA = 12'b010111100001;
            14'b10_000010110000: DATA = 12'b010111011110;
            14'b10_000010110001: DATA = 12'b010111011011;
            14'b10_000010110010: DATA = 12'b010111010111;
            14'b10_000010110011: DATA = 12'b010111010100;
            14'b10_000010110100: DATA = 12'b010111010001;
            14'b10_000010110101: DATA = 12'b010111001110;
            14'b10_000010110110: DATA = 12'b010111001011;
            14'b10_000010110111: DATA = 12'b010111001000;
            14'b10_000010111000: DATA = 12'b010111000101;
            14'b10_000010111001: DATA = 12'b010111000010;
            14'b10_000010111010: DATA = 12'b010110111111;
            14'b10_000010111011: DATA = 12'b010110111100;
            14'b10_000010111100: DATA = 12'b010110111001;
            14'b10_000010111101: DATA = 12'b010110110110;
            14'b10_000010111110: DATA = 12'b010110110011;
            14'b10_000010111111: DATA = 12'b010110110000;
            14'b10_000011000000: DATA = 12'b010110101101;
            14'b10_000011000001: DATA = 12'b010110101010;
            14'b10_000011000010: DATA = 12'b010110100111;
            14'b10_000011000011: DATA = 12'b010110100100;
            14'b10_000011000100: DATA = 12'b010110100001;
            14'b10_000011000101: DATA = 12'b010110011110;
            14'b10_000011000110: DATA = 12'b010110011011;
            14'b10_000011000111: DATA = 12'b010110011000;
            14'b10_000011001000: DATA = 12'b010110010101;
            14'b10_000011001001: DATA = 12'b010110010010;
            14'b10_000011001010: DATA = 12'b010110001111;
            14'b10_000011001011: DATA = 12'b010110001100;
            14'b10_000011001100: DATA = 12'b010110001001;
            14'b10_000011001101: DATA = 12'b010110000110;
            14'b10_000011001110: DATA = 12'b010110000011;
            14'b10_000011001111: DATA = 12'b010110000000;
            14'b10_000011010000: DATA = 12'b010101111101;
            14'b10_000011010001: DATA = 12'b010101111010;
            14'b10_000011010010: DATA = 12'b010101110111;
            14'b10_000011010011: DATA = 12'b010101110100;
            14'b10_000011010100: DATA = 12'b010101110001;
            14'b10_000011010101: DATA = 12'b010101101111;
            14'b10_000011010110: DATA = 12'b010101101100;
            14'b10_000011010111: DATA = 12'b010101101001;
            14'b10_000011011000: DATA = 12'b010101100110;
            14'b10_000011011001: DATA = 12'b010101100011;
            14'b10_000011011010: DATA = 12'b010101100000;
            14'b10_000011011011: DATA = 12'b010101011101;
            14'b10_000011011100: DATA = 12'b010101011010;
            14'b10_000011011101: DATA = 12'b010101010111;
            14'b10_000011011110: DATA = 12'b010101010100;
            14'b10_000011011111: DATA = 12'b010101010001;
            14'b10_000011100000: DATA = 12'b010101001110;
            14'b10_000011100001: DATA = 12'b010101001011;
            14'b10_000011100010: DATA = 12'b010101001000;
            14'b10_000011100011: DATA = 12'b010101000101;
            14'b10_000011100100: DATA = 12'b010101000010;
            14'b10_000011100101: DATA = 12'b010100111111;
            14'b10_000011100110: DATA = 12'b010100111100;
            14'b10_000011100111: DATA = 12'b010100111001;
            14'b10_000011101000: DATA = 12'b010100110110;
            14'b10_000011101001: DATA = 12'b010100110011;
            14'b10_000011101010: DATA = 12'b010100110000;
            14'b10_000011101011: DATA = 12'b010100101101;
            14'b10_000011101100: DATA = 12'b010100101011;
            14'b10_000011101101: DATA = 12'b010100101000;
            14'b10_000011101110: DATA = 12'b010100100101;
            14'b10_000011101111: DATA = 12'b010100100010;
            14'b10_000011110000: DATA = 12'b010100011111;
            14'b10_000011110001: DATA = 12'b010100011100;
            14'b10_000011110010: DATA = 12'b010100011001;
            14'b10_000011110011: DATA = 12'b010100010110;
            14'b10_000011110100: DATA = 12'b010100010011;
            14'b10_000011110101: DATA = 12'b010100010000;
            14'b10_000011110110: DATA = 12'b010100001101;
            14'b10_000011110111: DATA = 12'b010100001010;
            14'b10_000011111000: DATA = 12'b010100000111;
            14'b10_000011111001: DATA = 12'b010100000100;
            14'b10_000011111010: DATA = 12'b010100000010;
            14'b10_000011111011: DATA = 12'b010011111111;
            14'b10_000011111100: DATA = 12'b010011111100;
            14'b10_000011111101: DATA = 12'b010011111001;
            14'b10_000011111110: DATA = 12'b010011110110;
            14'b10_000011111111: DATA = 12'b010011110011;
            14'b10_000100000000: DATA = 12'b010011110000;
            14'b10_000100000001: DATA = 12'b010011101101;
            14'b10_000100000010: DATA = 12'b010011101010;
            14'b10_000100000011: DATA = 12'b010011100111;
            14'b10_000100000100: DATA = 12'b010011100101;
            14'b10_000100000101: DATA = 12'b010011100010;
            14'b10_000100000110: DATA = 12'b010011011111;
            14'b10_000100000111: DATA = 12'b010011011100;
            14'b10_000100001000: DATA = 12'b010011011001;
            14'b10_000100001001: DATA = 12'b010011010110;
            14'b10_000100001010: DATA = 12'b010011010011;
            14'b10_000100001011: DATA = 12'b010011010000;
            14'b10_000100001100: DATA = 12'b010011001101;
            14'b10_000100001101: DATA = 12'b010011001011;
            14'b10_000100001110: DATA = 12'b010011001000;
            14'b10_000100001111: DATA = 12'b010011000101;
            14'b10_000100010000: DATA = 12'b010011000010;
            14'b10_000100010001: DATA = 12'b010010111111;
            14'b10_000100010010: DATA = 12'b010010111100;
            14'b10_000100010011: DATA = 12'b010010111001;
            14'b10_000100010100: DATA = 12'b010010110111;
            14'b10_000100010101: DATA = 12'b010010110100;
            14'b10_000100010110: DATA = 12'b010010110001;
            14'b10_000100010111: DATA = 12'b010010101110;
            14'b10_000100011000: DATA = 12'b010010101011;
            14'b10_000100011001: DATA = 12'b010010101000;
            14'b10_000100011010: DATA = 12'b010010100101;
            14'b10_000100011011: DATA = 12'b010010100011;
            14'b10_000100011100: DATA = 12'b010010100000;
            14'b10_000100011101: DATA = 12'b010010011101;
            14'b10_000100011110: DATA = 12'b010010011010;
            14'b10_000100011111: DATA = 12'b010010010111;
            14'b10_000100100000: DATA = 12'b010010010100;
            14'b10_000100100001: DATA = 12'b010010010001;
            14'b10_000100100010: DATA = 12'b010010001111;
            14'b10_000100100011: DATA = 12'b010010001100;
            14'b10_000100100100: DATA = 12'b010010001001;
            14'b10_000100100101: DATA = 12'b010010000110;
            14'b10_000100100110: DATA = 12'b010010000011;
            14'b10_000100100111: DATA = 12'b010010000000;
            14'b10_000100101000: DATA = 12'b010001111110;
            14'b10_000100101001: DATA = 12'b010001111011;
            14'b10_000100101010: DATA = 12'b010001111000;
            14'b10_000100101011: DATA = 12'b010001110101;
            14'b10_000100101100: DATA = 12'b010001110010;
            14'b10_000100101101: DATA = 12'b010001110000;
            14'b10_000100101110: DATA = 12'b010001101101;
            14'b10_000100101111: DATA = 12'b010001101010;
            14'b10_000100110000: DATA = 12'b010001100111;
            14'b10_000100110001: DATA = 12'b010001100100;
            14'b10_000100110010: DATA = 12'b010001100010;
            14'b10_000100110011: DATA = 12'b010001011111;
            14'b10_000100110100: DATA = 12'b010001011100;
            14'b10_000100110101: DATA = 12'b010001011001;
            14'b10_000100110110: DATA = 12'b010001010110;
            14'b10_000100110111: DATA = 12'b010001010100;
            14'b10_000100111000: DATA = 12'b010001010001;
            14'b10_000100111001: DATA = 12'b010001001110;
            14'b10_000100111010: DATA = 12'b010001001011;
            14'b10_000100111011: DATA = 12'b010001001000;
            14'b10_000100111100: DATA = 12'b010001000110;
            14'b10_000100111101: DATA = 12'b010001000011;
            14'b10_000100111110: DATA = 12'b010001000000;
            14'b10_000100111111: DATA = 12'b010000111101;
            14'b10_000101000000: DATA = 12'b010000111011;
            14'b10_000101000001: DATA = 12'b010000111000;
            14'b10_000101000010: DATA = 12'b010000110101;
            14'b10_000101000011: DATA = 12'b010000110010;
            14'b10_000101000100: DATA = 12'b010000101111;
            14'b10_000101000101: DATA = 12'b010000101101;
            14'b10_000101000110: DATA = 12'b010000101010;
            14'b10_000101000111: DATA = 12'b010000100111;
            14'b10_000101001000: DATA = 12'b010000100100;
            14'b10_000101001001: DATA = 12'b010000100010;
            14'b10_000101001010: DATA = 12'b010000011111;
            14'b10_000101001011: DATA = 12'b010000011100;
            14'b10_000101001100: DATA = 12'b010000011001;
            14'b10_000101001101: DATA = 12'b010000010111;
            14'b10_000101001110: DATA = 12'b010000010100;
            14'b10_000101001111: DATA = 12'b010000010001;
            14'b10_000101010000: DATA = 12'b010000001111;
            14'b10_000101010001: DATA = 12'b010000001100;
            14'b10_000101010010: DATA = 12'b010000001001;
            14'b10_000101010011: DATA = 12'b010000000110;
            14'b10_000101010100: DATA = 12'b010000000100;
            14'b10_000101010101: DATA = 12'b010000000001;
            14'b10_000101010110: DATA = 12'b001111111110;
            14'b10_000101010111: DATA = 12'b001111111011;
            14'b10_000101011000: DATA = 12'b001111111001;
            14'b10_000101011001: DATA = 12'b001111110110;
            14'b10_000101011010: DATA = 12'b001111110011;
            14'b10_000101011011: DATA = 12'b001111110001;
            14'b10_000101011100: DATA = 12'b001111101110;
            14'b10_000101011101: DATA = 12'b001111101011;
            14'b10_000101011110: DATA = 12'b001111101001;
            14'b10_000101011111: DATA = 12'b001111100110;
            14'b10_000101100000: DATA = 12'b001111100011;
            14'b10_000101100001: DATA = 12'b001111100000;
            14'b10_000101100010: DATA = 12'b001111011110;
            14'b10_000101100011: DATA = 12'b001111011011;
            14'b10_000101100100: DATA = 12'b001111011000;
            14'b10_000101100101: DATA = 12'b001111010110;
            14'b10_000101100110: DATA = 12'b001111010011;
            14'b10_000101100111: DATA = 12'b001111010000;
            14'b10_000101101000: DATA = 12'b001111001110;
            14'b10_000101101001: DATA = 12'b001111001011;
            14'b10_000101101010: DATA = 12'b001111001000;
            14'b10_000101101011: DATA = 12'b001111000110;
            14'b10_000101101100: DATA = 12'b001111000011;
            14'b10_000101101101: DATA = 12'b001111000000;
            14'b10_000101101110: DATA = 12'b001110111110;
            14'b10_000101101111: DATA = 12'b001110111011;
            14'b10_000101110000: DATA = 12'b001110111000;
            14'b10_000101110001: DATA = 12'b001110110110;
            14'b10_000101110010: DATA = 12'b001110110011;
            14'b10_000101110011: DATA = 12'b001110110000;
            14'b10_000101110100: DATA = 12'b001110101110;
            14'b10_000101110101: DATA = 12'b001110101011;
            14'b10_000101110110: DATA = 12'b001110101000;
            14'b10_000101110111: DATA = 12'b001110100110;
            14'b10_000101111000: DATA = 12'b001110100011;
            14'b10_000101111001: DATA = 12'b001110100001;
            14'b10_000101111010: DATA = 12'b001110011110;
            14'b10_000101111011: DATA = 12'b001110011011;
            14'b10_000101111100: DATA = 12'b001110011001;
            14'b10_000101111101: DATA = 12'b001110010110;
            14'b10_000101111110: DATA = 12'b001110010011;
            14'b10_000101111111: DATA = 12'b001110010001;
            14'b10_000110000000: DATA = 12'b001110001110;
            14'b10_000110000001: DATA = 12'b001110001100;
            14'b10_000110000010: DATA = 12'b001110001001;
            14'b10_000110000011: DATA = 12'b001110000110;
            14'b10_000110000100: DATA = 12'b001110000100;
            14'b10_000110000101: DATA = 12'b001110000001;
            14'b10_000110000110: DATA = 12'b001101111111;
            14'b10_000110000111: DATA = 12'b001101111100;
            14'b10_000110001000: DATA = 12'b001101111001;
            14'b10_000110001001: DATA = 12'b001101110111;
            14'b10_000110001010: DATA = 12'b001101110100;
            14'b10_000110001011: DATA = 12'b001101110010;
            14'b10_000110001100: DATA = 12'b001101101111;
            14'b10_000110001101: DATA = 12'b001101101101;
            14'b10_000110001110: DATA = 12'b001101101010;
            14'b10_000110001111: DATA = 12'b001101100111;
            14'b10_000110010000: DATA = 12'b001101100101;
            14'b10_000110010001: DATA = 12'b001101100010;
            14'b10_000110010010: DATA = 12'b001101100000;
            14'b10_000110010011: DATA = 12'b001101011101;
            14'b10_000110010100: DATA = 12'b001101011011;
            14'b10_000110010101: DATA = 12'b001101011000;
            14'b10_000110010110: DATA = 12'b001101010101;
            14'b10_000110010111: DATA = 12'b001101010011;
            14'b10_000110011000: DATA = 12'b001101010000;
            14'b10_000110011001: DATA = 12'b001101001110;
            14'b10_000110011010: DATA = 12'b001101001011;
            14'b10_000110011011: DATA = 12'b001101001001;
            14'b10_000110011100: DATA = 12'b001101000110;
            14'b10_000110011101: DATA = 12'b001101000100;
            14'b10_000110011110: DATA = 12'b001101000001;
            14'b10_000110011111: DATA = 12'b001100111111;
            14'b10_000110100000: DATA = 12'b001100111100;
            14'b10_000110100001: DATA = 12'b001100111010;
            14'b10_000110100010: DATA = 12'b001100110111;
            14'b10_000110100011: DATA = 12'b001100110101;
            14'b10_000110100100: DATA = 12'b001100110010;
            14'b10_000110100101: DATA = 12'b001100110000;
            14'b10_000110100110: DATA = 12'b001100101101;
            14'b10_000110100111: DATA = 12'b001100101011;
            14'b10_000110101000: DATA = 12'b001100101000;
            14'b10_000110101001: DATA = 12'b001100100110;
            14'b10_000110101010: DATA = 12'b001100100011;
            14'b10_000110101011: DATA = 12'b001100100001;
            14'b10_000110101100: DATA = 12'b001100011110;
            14'b10_000110101101: DATA = 12'b001100011100;
            14'b10_000110101110: DATA = 12'b001100011001;
            14'b10_000110101111: DATA = 12'b001100010111;
            14'b10_000110110000: DATA = 12'b001100010100;
            14'b10_000110110001: DATA = 12'b001100010010;
            14'b10_000110110010: DATA = 12'b001100001111;
            14'b10_000110110011: DATA = 12'b001100001101;
            14'b10_000110110100: DATA = 12'b001100001010;
            14'b10_000110110101: DATA = 12'b001100001000;
            14'b10_000110110110: DATA = 12'b001100000101;
            14'b10_000110110111: DATA = 12'b001100000011;
            14'b10_000110111000: DATA = 12'b001100000000;
            14'b10_000110111001: DATA = 12'b001011111110;
            14'b10_000110111010: DATA = 12'b001011111100;
            14'b10_000110111011: DATA = 12'b001011111001;
            14'b10_000110111100: DATA = 12'b001011110111;
            14'b10_000110111101: DATA = 12'b001011110100;
            14'b10_000110111110: DATA = 12'b001011110010;
            14'b10_000110111111: DATA = 12'b001011101111;
            14'b10_000111000000: DATA = 12'b001011101101;
            14'b10_000111000001: DATA = 12'b001011101010;
            14'b10_000111000010: DATA = 12'b001011101000;
            14'b10_000111000011: DATA = 12'b001011100110;
            14'b10_000111000100: DATA = 12'b001011100011;
            14'b10_000111000101: DATA = 12'b001011100001;
            14'b10_000111000110: DATA = 12'b001011011110;
            14'b10_000111000111: DATA = 12'b001011011100;
            14'b10_000111001000: DATA = 12'b001011011010;
            14'b10_000111001001: DATA = 12'b001011010111;
            14'b10_000111001010: DATA = 12'b001011010101;
            14'b10_000111001011: DATA = 12'b001011010010;
            14'b10_000111001100: DATA = 12'b001011010000;
            14'b10_000111001101: DATA = 12'b001011001110;
            14'b10_000111001110: DATA = 12'b001011001011;
            14'b10_000111001111: DATA = 12'b001011001001;
            14'b10_000111010000: DATA = 12'b001011000110;
            14'b10_000111010001: DATA = 12'b001011000100;
            14'b10_000111010010: DATA = 12'b001011000010;
            14'b10_000111010011: DATA = 12'b001010111111;
            14'b10_000111010100: DATA = 12'b001010111101;
            14'b10_000111010101: DATA = 12'b001010111011;
            14'b10_000111010110: DATA = 12'b001010111000;
            14'b10_000111010111: DATA = 12'b001010110110;
            14'b10_000111011000: DATA = 12'b001010110100;
            14'b10_000111011001: DATA = 12'b001010110001;
            14'b10_000111011010: DATA = 12'b001010101111;
            14'b10_000111011011: DATA = 12'b001010101100;
            14'b10_000111011100: DATA = 12'b001010101010;
            14'b10_000111011101: DATA = 12'b001010101000;
            14'b10_000111011110: DATA = 12'b001010100101;
            14'b10_000111011111: DATA = 12'b001010100011;
            14'b10_000111100000: DATA = 12'b001010100001;
            14'b10_000111100001: DATA = 12'b001010011110;
            14'b10_000111100010: DATA = 12'b001010011100;
            14'b10_000111100011: DATA = 12'b001010011010;
            14'b10_000111100100: DATA = 12'b001010011000;
            14'b10_000111100101: DATA = 12'b001010010101;
            14'b10_000111100110: DATA = 12'b001010010011;
            14'b10_000111100111: DATA = 12'b001010010001;
            14'b10_000111101000: DATA = 12'b001010001110;
            14'b10_000111101001: DATA = 12'b001010001100;
            14'b10_000111101010: DATA = 12'b001010001010;
            14'b10_000111101011: DATA = 12'b001010000111;
            14'b10_000111101100: DATA = 12'b001010000101;
            14'b10_000111101101: DATA = 12'b001010000011;
            14'b10_000111101110: DATA = 12'b001010000001;
            14'b10_000111101111: DATA = 12'b001001111110;
            14'b10_000111110000: DATA = 12'b001001111100;
            14'b10_000111110001: DATA = 12'b001001111010;
            14'b10_000111110010: DATA = 12'b001001110111;
            14'b10_000111110011: DATA = 12'b001001110101;
            14'b10_000111110100: DATA = 12'b001001110011;
            14'b10_000111110101: DATA = 12'b001001110001;
            14'b10_000111110110: DATA = 12'b001001101110;
            14'b10_000111110111: DATA = 12'b001001101100;
            14'b10_000111111000: DATA = 12'b001001101010;
            14'b10_000111111001: DATA = 12'b001001101000;
            14'b10_000111111010: DATA = 12'b001001100101;
            14'b10_000111111011: DATA = 12'b001001100011;
            14'b10_000111111100: DATA = 12'b001001100001;
            14'b10_000111111101: DATA = 12'b001001011111;
            14'b10_000111111110: DATA = 12'b001001011100;
            14'b10_000111111111: DATA = 12'b001001011010;
            14'b10_001000000000: DATA = 12'b001001011000;
            14'b10_001000000001: DATA = 12'b001001010110;
            14'b10_001000000010: DATA = 12'b001001010100;
            14'b10_001000000011: DATA = 12'b001001010001;
            14'b10_001000000100: DATA = 12'b001001001111;
            14'b10_001000000101: DATA = 12'b001001001101;
            14'b10_001000000110: DATA = 12'b001001001011;
            14'b10_001000000111: DATA = 12'b001001001001;
            14'b10_001000001000: DATA = 12'b001001000110;
            14'b10_001000001001: DATA = 12'b001001000100;
            14'b10_001000001010: DATA = 12'b001001000010;
            14'b10_001000001011: DATA = 12'b001001000000;
            14'b10_001000001100: DATA = 12'b001000111110;
            14'b10_001000001101: DATA = 12'b001000111011;
            14'b10_001000001110: DATA = 12'b001000111001;
            14'b10_001000001111: DATA = 12'b001000110111;
            14'b10_001000010000: DATA = 12'b001000110101;
            14'b10_001000010001: DATA = 12'b001000110011;
            14'b10_001000010010: DATA = 12'b001000110001;
            14'b10_001000010011: DATA = 12'b001000101110;
            14'b10_001000010100: DATA = 12'b001000101100;
            14'b10_001000010101: DATA = 12'b001000101010;
            14'b10_001000010110: DATA = 12'b001000101000;
            14'b10_001000010111: DATA = 12'b001000100110;
            14'b10_001000011000: DATA = 12'b001000100100;
            14'b10_001000011001: DATA = 12'b001000100010;
            14'b10_001000011010: DATA = 12'b001000011111;
            14'b10_001000011011: DATA = 12'b001000011101;
            14'b10_001000011100: DATA = 12'b001000011011;
            14'b10_001000011101: DATA = 12'b001000011001;
            14'b10_001000011110: DATA = 12'b001000010111;
            14'b10_001000011111: DATA = 12'b001000010101;
            14'b10_001000100000: DATA = 12'b001000010011;
            14'b10_001000100001: DATA = 12'b001000010001;
            14'b10_001000100010: DATA = 12'b001000001111;
            14'b10_001000100011: DATA = 12'b001000001100;
            14'b10_001000100100: DATA = 12'b001000001010;
            14'b10_001000100101: DATA = 12'b001000001000;
            14'b10_001000100110: DATA = 12'b001000000110;
            14'b10_001000100111: DATA = 12'b001000000100;
            14'b10_001000101000: DATA = 12'b001000000010;
            14'b10_001000101001: DATA = 12'b001000000000;
            14'b10_001000101010: DATA = 12'b000111111110;
            14'b10_001000101011: DATA = 12'b000111111100;
            14'b10_001000101100: DATA = 12'b000111111010;
            14'b10_001000101101: DATA = 12'b000111111000;
            14'b10_001000101110: DATA = 12'b000111110110;
            14'b10_001000101111: DATA = 12'b000111110100;
            14'b10_001000110000: DATA = 12'b000111110001;
            14'b10_001000110001: DATA = 12'b000111101111;
            14'b10_001000110010: DATA = 12'b000111101101;
            14'b10_001000110011: DATA = 12'b000111101011;
            14'b10_001000110100: DATA = 12'b000111101001;
            14'b10_001000110101: DATA = 12'b000111100111;
            14'b10_001000110110: DATA = 12'b000111100101;
            14'b10_001000110111: DATA = 12'b000111100011;
            14'b10_001000111000: DATA = 12'b000111100001;
            14'b10_001000111001: DATA = 12'b000111011111;
            14'b10_001000111010: DATA = 12'b000111011101;
            14'b10_001000111011: DATA = 12'b000111011011;
            14'b10_001000111100: DATA = 12'b000111011001;
            14'b10_001000111101: DATA = 12'b000111010111;
            14'b10_001000111110: DATA = 12'b000111010101;
            14'b10_001000111111: DATA = 12'b000111010011;
            14'b10_001001000000: DATA = 12'b000111010001;
            14'b10_001001000001: DATA = 12'b000111001111;
            14'b10_001001000010: DATA = 12'b000111001101;
            14'b10_001001000011: DATA = 12'b000111001011;
            14'b10_001001000100: DATA = 12'b000111001001;
            14'b10_001001000101: DATA = 12'b000111000111;
            14'b10_001001000110: DATA = 12'b000111000101;
            14'b10_001001000111: DATA = 12'b000111000011;
            14'b10_001001001000: DATA = 12'b000111000001;
            14'b10_001001001001: DATA = 12'b000110111111;
            14'b10_001001001010: DATA = 12'b000110111101;
            14'b10_001001001011: DATA = 12'b000110111011;
            14'b10_001001001100: DATA = 12'b000110111010;
            14'b10_001001001101: DATA = 12'b000110111000;
            14'b10_001001001110: DATA = 12'b000110110110;
            14'b10_001001001111: DATA = 12'b000110110100;
            14'b10_001001010000: DATA = 12'b000110110010;
            14'b10_001001010001: DATA = 12'b000110110000;
            14'b10_001001010010: DATA = 12'b000110101110;
            14'b10_001001010011: DATA = 12'b000110101100;
            14'b10_001001010100: DATA = 12'b000110101010;
            14'b10_001001010101: DATA = 12'b000110101000;
            14'b10_001001010110: DATA = 12'b000110100110;
            14'b10_001001010111: DATA = 12'b000110100100;
            14'b10_001001011000: DATA = 12'b000110100010;
            14'b10_001001011001: DATA = 12'b000110100001;
            14'b10_001001011010: DATA = 12'b000110011111;
            14'b10_001001011011: DATA = 12'b000110011101;
            14'b10_001001011100: DATA = 12'b000110011011;
            14'b10_001001011101: DATA = 12'b000110011001;
            14'b10_001001011110: DATA = 12'b000110010111;
            14'b10_001001011111: DATA = 12'b000110010101;
            14'b10_001001100000: DATA = 12'b000110010011;
            14'b10_001001100001: DATA = 12'b000110010001;
            14'b10_001001100010: DATA = 12'b000110010000;
            14'b10_001001100011: DATA = 12'b000110001110;
            14'b10_001001100100: DATA = 12'b000110001100;
            14'b10_001001100101: DATA = 12'b000110001010;
            14'b10_001001100110: DATA = 12'b000110001000;
            14'b10_001001100111: DATA = 12'b000110000110;
            14'b10_001001101000: DATA = 12'b000110000100;
            14'b10_001001101001: DATA = 12'b000110000011;
            14'b10_001001101010: DATA = 12'b000110000001;
            14'b10_001001101011: DATA = 12'b000101111111;
            14'b10_001001101100: DATA = 12'b000101111101;
            14'b10_001001101101: DATA = 12'b000101111011;
            14'b10_001001101110: DATA = 12'b000101111010;
            14'b10_001001101111: DATA = 12'b000101111000;
            14'b10_001001110000: DATA = 12'b000101110110;
            14'b10_001001110001: DATA = 12'b000101110100;
            14'b10_001001110010: DATA = 12'b000101110010;
            14'b10_001001110011: DATA = 12'b000101110000;
            14'b10_001001110100: DATA = 12'b000101101111;
            14'b10_001001110101: DATA = 12'b000101101101;
            14'b10_001001110110: DATA = 12'b000101101011;
            14'b10_001001110111: DATA = 12'b000101101001;
            14'b10_001001111000: DATA = 12'b000101101000;
            14'b10_001001111001: DATA = 12'b000101100110;
            14'b10_001001111010: DATA = 12'b000101100100;
            14'b10_001001111011: DATA = 12'b000101100010;
            14'b10_001001111100: DATA = 12'b000101100000;
            14'b10_001001111101: DATA = 12'b000101011111;
            14'b10_001001111110: DATA = 12'b000101011101;
            14'b10_001001111111: DATA = 12'b000101011011;
            14'b10_001010000000: DATA = 12'b000101011001;
            14'b10_001010000001: DATA = 12'b000101011000;
            14'b10_001010000010: DATA = 12'b000101010110;
            14'b10_001010000011: DATA = 12'b000101010100;
            14'b10_001010000100: DATA = 12'b000101010011;
            14'b10_001010000101: DATA = 12'b000101010001;
            14'b10_001010000110: DATA = 12'b000101001111;
            14'b10_001010000111: DATA = 12'b000101001101;
            14'b10_001010001000: DATA = 12'b000101001100;
            14'b10_001010001001: DATA = 12'b000101001010;
            14'b10_001010001010: DATA = 12'b000101001000;
            14'b10_001010001011: DATA = 12'b000101000111;
            14'b10_001010001100: DATA = 12'b000101000101;
            14'b10_001010001101: DATA = 12'b000101000011;
            14'b10_001010001110: DATA = 12'b000101000001;
            14'b10_001010001111: DATA = 12'b000101000000;
            14'b10_001010010000: DATA = 12'b000100111110;
            14'b10_001010010001: DATA = 12'b000100111100;
            14'b10_001010010010: DATA = 12'b000100111011;
            14'b10_001010010011: DATA = 12'b000100111001;
            14'b10_001010010100: DATA = 12'b000100110111;
            14'b10_001010010101: DATA = 12'b000100110110;
            14'b10_001010010110: DATA = 12'b000100110100;
            14'b10_001010010111: DATA = 12'b000100110010;
            14'b10_001010011000: DATA = 12'b000100110001;
            14'b10_001010011001: DATA = 12'b000100101111;
            14'b10_001010011010: DATA = 12'b000100101101;
            14'b10_001010011011: DATA = 12'b000100101100;
            14'b10_001010011100: DATA = 12'b000100101010;
            14'b10_001010011101: DATA = 12'b000100101001;
            14'b10_001010011110: DATA = 12'b000100100111;
            14'b10_001010011111: DATA = 12'b000100100101;
            14'b10_001010100000: DATA = 12'b000100100100;
            14'b10_001010100001: DATA = 12'b000100100010;
            14'b10_001010100010: DATA = 12'b000100100001;
            14'b10_001010100011: DATA = 12'b000100011111;
            14'b10_001010100100: DATA = 12'b000100011101;
            14'b10_001010100101: DATA = 12'b000100011100;
            14'b10_001010100110: DATA = 12'b000100011010;
            14'b10_001010100111: DATA = 12'b000100011001;
            14'b10_001010101000: DATA = 12'b000100010111;
            14'b10_001010101001: DATA = 12'b000100010101;
            14'b10_001010101010: DATA = 12'b000100010100;
            14'b10_001010101011: DATA = 12'b000100010010;
            14'b10_001010101100: DATA = 12'b000100010001;
            14'b10_001010101101: DATA = 12'b000100001111;
            14'b10_001010101110: DATA = 12'b000100001110;
            14'b10_001010101111: DATA = 12'b000100001100;
            14'b10_001010110000: DATA = 12'b000100001010;
            14'b10_001010110001: DATA = 12'b000100001001;
            14'b10_001010110010: DATA = 12'b000100000111;
            14'b10_001010110011: DATA = 12'b000100000110;
            14'b10_001010110100: DATA = 12'b000100000100;
            14'b10_001010110101: DATA = 12'b000100000011;
            14'b10_001010110110: DATA = 12'b000100000001;
            14'b10_001010110111: DATA = 12'b000100000000;
            14'b10_001010111000: DATA = 12'b000011111110;
            14'b10_001010111001: DATA = 12'b000011111101;
            14'b10_001010111010: DATA = 12'b000011111011;
            14'b10_001010111011: DATA = 12'b000011111010;
            14'b10_001010111100: DATA = 12'b000011111000;
            14'b10_001010111101: DATA = 12'b000011110111;
            14'b10_001010111110: DATA = 12'b000011110101;
            14'b10_001010111111: DATA = 12'b000011110100;
            14'b10_001011000000: DATA = 12'b000011110010;
            14'b10_001011000001: DATA = 12'b000011110001;
            14'b10_001011000010: DATA = 12'b000011101111;
            14'b10_001011000011: DATA = 12'b000011101110;
            14'b10_001011000100: DATA = 12'b000011101100;
            14'b10_001011000101: DATA = 12'b000011101011;
            14'b10_001011000110: DATA = 12'b000011101001;
            14'b10_001011000111: DATA = 12'b000011101000;
            14'b10_001011001000: DATA = 12'b000011100111;
            14'b10_001011001001: DATA = 12'b000011100101;
            14'b10_001011001010: DATA = 12'b000011100100;
            14'b10_001011001011: DATA = 12'b000011100010;
            14'b10_001011001100: DATA = 12'b000011100001;
            14'b10_001011001101: DATA = 12'b000011011111;
            14'b10_001011001110: DATA = 12'b000011011110;
            14'b10_001011001111: DATA = 12'b000011011100;
            14'b10_001011010000: DATA = 12'b000011011011;
            14'b10_001011010001: DATA = 12'b000011011010;
            14'b10_001011010010: DATA = 12'b000011011000;
            14'b10_001011010011: DATA = 12'b000011010111;
            14'b10_001011010100: DATA = 12'b000011010101;
            14'b10_001011010101: DATA = 12'b000011010100;
            14'b10_001011010110: DATA = 12'b000011010011;
            14'b10_001011010111: DATA = 12'b000011010001;
            14'b10_001011011000: DATA = 12'b000011010000;
            14'b10_001011011001: DATA = 12'b000011001111;
            14'b10_001011011010: DATA = 12'b000011001101;
            14'b10_001011011011: DATA = 12'b000011001100;
            14'b10_001011011100: DATA = 12'b000011001010;
            14'b10_001011011101: DATA = 12'b000011001001;
            14'b10_001011011110: DATA = 12'b000011001000;
            14'b10_001011011111: DATA = 12'b000011000110;
            14'b10_001011100000: DATA = 12'b000011000101;
            14'b10_001011100001: DATA = 12'b000011000100;
            14'b10_001011100010: DATA = 12'b000011000010;
            14'b10_001011100011: DATA = 12'b000011000001;
            14'b10_001011100100: DATA = 12'b000011000000;
            14'b10_001011100101: DATA = 12'b000010111110;
            14'b10_001011100110: DATA = 12'b000010111101;
            14'b10_001011100111: DATA = 12'b000010111100;
            14'b10_001011101000: DATA = 12'b000010111010;
            14'b10_001011101001: DATA = 12'b000010111001;
            14'b10_001011101010: DATA = 12'b000010111000;
            14'b10_001011101011: DATA = 12'b000010110111;
            14'b10_001011101100: DATA = 12'b000010110101;
            14'b10_001011101101: DATA = 12'b000010110100;
            14'b10_001011101110: DATA = 12'b000010110011;
            14'b10_001011101111: DATA = 12'b000010110001;
            14'b10_001011110000: DATA = 12'b000010110000;
            14'b10_001011110001: DATA = 12'b000010101111;
            14'b10_001011110010: DATA = 12'b000010101110;
            14'b10_001011110011: DATA = 12'b000010101100;
            14'b10_001011110100: DATA = 12'b000010101011;
            14'b10_001011110101: DATA = 12'b000010101010;
            14'b10_001011110110: DATA = 12'b000010101001;
            14'b10_001011110111: DATA = 12'b000010100111;
            14'b10_001011111000: DATA = 12'b000010100110;
            14'b10_001011111001: DATA = 12'b000010100101;
            14'b10_001011111010: DATA = 12'b000010100100;
            14'b10_001011111011: DATA = 12'b000010100010;
            14'b10_001011111100: DATA = 12'b000010100001;
            14'b10_001011111101: DATA = 12'b000010100000;
            14'b10_001011111110: DATA = 12'b000010011111;
            14'b10_001011111111: DATA = 12'b000010011110;
            14'b10_001100000000: DATA = 12'b000010011100;
            14'b10_001100000001: DATA = 12'b000010011011;
            14'b10_001100000010: DATA = 12'b000010011010;
            14'b10_001100000011: DATA = 12'b000010011001;
            14'b10_001100000100: DATA = 12'b000010011000;
            14'b10_001100000101: DATA = 12'b000010010110;
            14'b10_001100000110: DATA = 12'b000010010101;
            14'b10_001100000111: DATA = 12'b000010010100;
            14'b10_001100001000: DATA = 12'b000010010011;
            14'b10_001100001001: DATA = 12'b000010010010;
            14'b10_001100001010: DATA = 12'b000010010001;
            14'b10_001100001011: DATA = 12'b000010001111;
            14'b10_001100001100: DATA = 12'b000010001110;
            14'b10_001100001101: DATA = 12'b000010001101;
            14'b10_001100001110: DATA = 12'b000010001100;
            14'b10_001100001111: DATA = 12'b000010001011;
            14'b10_001100010000: DATA = 12'b000010001010;
            14'b10_001100010001: DATA = 12'b000010001001;
            14'b10_001100010010: DATA = 12'b000010000111;
            14'b10_001100010011: DATA = 12'b000010000110;
            14'b10_001100010100: DATA = 12'b000010000101;
            14'b10_001100010101: DATA = 12'b000010000100;
            14'b10_001100010110: DATA = 12'b000010000011;
            14'b10_001100010111: DATA = 12'b000010000010;
            14'b10_001100011000: DATA = 12'b000010000001;
            14'b10_001100011001: DATA = 12'b000010000000;
            14'b10_001100011010: DATA = 12'b000001111111;
            14'b10_001100011011: DATA = 12'b000001111110;
            14'b10_001100011100: DATA = 12'b000001111100;
            14'b10_001100011101: DATA = 12'b000001111011;
            14'b10_001100011110: DATA = 12'b000001111010;
            14'b10_001100011111: DATA = 12'b000001111001;
            14'b10_001100100000: DATA = 12'b000001111000;
            14'b10_001100100001: DATA = 12'b000001110111;
            14'b10_001100100010: DATA = 12'b000001110110;
            14'b10_001100100011: DATA = 12'b000001110101;
            14'b10_001100100100: DATA = 12'b000001110100;
            14'b10_001100100101: DATA = 12'b000001110011;
            14'b10_001100100110: DATA = 12'b000001110010;
            14'b10_001100100111: DATA = 12'b000001110001;
            14'b10_001100101000: DATA = 12'b000001110000;
            14'b10_001100101001: DATA = 12'b000001101111;
            14'b10_001100101010: DATA = 12'b000001101110;
            14'b10_001100101011: DATA = 12'b000001101101;
            14'b10_001100101100: DATA = 12'b000001101100;
            14'b10_001100101101: DATA = 12'b000001101011;
            14'b10_001100101110: DATA = 12'b000001101010;
            14'b10_001100101111: DATA = 12'b000001101001;
            14'b10_001100110000: DATA = 12'b000001101000;
            14'b10_001100110001: DATA = 12'b000001100111;
            14'b10_001100110010: DATA = 12'b000001100110;
            14'b10_001100110011: DATA = 12'b000001100101;
            14'b10_001100110100: DATA = 12'b000001100100;
            14'b10_001100110101: DATA = 12'b000001100011;
            14'b10_001100110110: DATA = 12'b000001100010;
            14'b10_001100110111: DATA = 12'b000001100001;
            14'b10_001100111000: DATA = 12'b000001100000;
            14'b10_001100111001: DATA = 12'b000001011111;
            14'b10_001100111010: DATA = 12'b000001011110;
            14'b10_001100111011: DATA = 12'b000001011101;
            14'b10_001100111100: DATA = 12'b000001011100;
            14'b10_001100111101: DATA = 12'b000001011011;
            14'b10_001100111110: DATA = 12'b000001011010;
            14'b10_001100111111: DATA = 12'b000001011010;
            14'b10_001101000000: DATA = 12'b000001011001;
            14'b10_001101000001: DATA = 12'b000001011000;
            14'b10_001101000010: DATA = 12'b000001010111;
            14'b10_001101000011: DATA = 12'b000001010110;
            14'b10_001101000100: DATA = 12'b000001010101;
            14'b10_001101000101: DATA = 12'b000001010100;
            14'b10_001101000110: DATA = 12'b000001010011;
            14'b10_001101000111: DATA = 12'b000001010010;
            14'b10_001101001000: DATA = 12'b000001010001;
            14'b10_001101001001: DATA = 12'b000001010001;
            14'b10_001101001010: DATA = 12'b000001010000;
            14'b10_001101001011: DATA = 12'b000001001111;
            14'b10_001101001100: DATA = 12'b000001001110;
            14'b10_001101001101: DATA = 12'b000001001101;
            14'b10_001101001110: DATA = 12'b000001001100;
            14'b10_001101001111: DATA = 12'b000001001011;
            14'b10_001101010000: DATA = 12'b000001001011;
            14'b10_001101010001: DATA = 12'b000001001010;
            14'b10_001101010010: DATA = 12'b000001001001;
            14'b10_001101010011: DATA = 12'b000001001000;
            14'b10_001101010100: DATA = 12'b000001000111;
            14'b10_001101010101: DATA = 12'b000001000111;
            14'b10_001101010110: DATA = 12'b000001000110;
            14'b10_001101010111: DATA = 12'b000001000101;
            14'b10_001101011000: DATA = 12'b000001000100;
            14'b10_001101011001: DATA = 12'b000001000011;
            14'b10_001101011010: DATA = 12'b000001000011;
            14'b10_001101011011: DATA = 12'b000001000010;
            14'b10_001101011100: DATA = 12'b000001000001;
            14'b10_001101011101: DATA = 12'b000001000000;
            14'b10_001101011110: DATA = 12'b000000111111;
            14'b10_001101011111: DATA = 12'b000000111111;
            14'b10_001101100000: DATA = 12'b000000111110;
            14'b10_001101100001: DATA = 12'b000000111101;
            14'b10_001101100010: DATA = 12'b000000111100;
            14'b10_001101100011: DATA = 12'b000000111100;
            14'b10_001101100100: DATA = 12'b000000111011;
            14'b10_001101100101: DATA = 12'b000000111010;
            14'b10_001101100110: DATA = 12'b000000111001;
            14'b10_001101100111: DATA = 12'b000000111001;
            14'b10_001101101000: DATA = 12'b000000111000;
            14'b10_001101101001: DATA = 12'b000000110111;
            14'b10_001101101010: DATA = 12'b000000110110;
            14'b10_001101101011: DATA = 12'b000000110110;
            14'b10_001101101100: DATA = 12'b000000110101;
            14'b10_001101101101: DATA = 12'b000000110100;
            14'b10_001101101110: DATA = 12'b000000110100;
            14'b10_001101101111: DATA = 12'b000000110011;
            14'b10_001101110000: DATA = 12'b000000110010;
            14'b10_001101110001: DATA = 12'b000000110010;
            14'b10_001101110010: DATA = 12'b000000110001;
            14'b10_001101110011: DATA = 12'b000000110000;
            14'b10_001101110100: DATA = 12'b000000110000;
            14'b10_001101110101: DATA = 12'b000000101111;
            14'b10_001101110110: DATA = 12'b000000101110;
            14'b10_001101110111: DATA = 12'b000000101110;
            14'b10_001101111000: DATA = 12'b000000101101;
            14'b10_001101111001: DATA = 12'b000000101100;
            14'b10_001101111010: DATA = 12'b000000101100;
            14'b10_001101111011: DATA = 12'b000000101011;
            14'b10_001101111100: DATA = 12'b000000101010;
            14'b10_001101111101: DATA = 12'b000000101010;
            14'b10_001101111110: DATA = 12'b000000101001;
            14'b10_001101111111: DATA = 12'b000000101000;
            14'b10_001110000000: DATA = 12'b000000101000;
            14'b10_001110000001: DATA = 12'b000000100111;
            14'b10_001110000010: DATA = 12'b000000100111;
            14'b10_001110000011: DATA = 12'b000000100110;
            14'b10_001110000100: DATA = 12'b000000100101;
            14'b10_001110000101: DATA = 12'b000000100101;
            14'b10_001110000110: DATA = 12'b000000100100;
            14'b10_001110000111: DATA = 12'b000000100100;
            14'b10_001110001000: DATA = 12'b000000100011;
            14'b10_001110001001: DATA = 12'b000000100011;
            14'b10_001110001010: DATA = 12'b000000100010;
            14'b10_001110001011: DATA = 12'b000000100001;
            14'b10_001110001100: DATA = 12'b000000100001;
            14'b10_001110001101: DATA = 12'b000000100000;
            14'b10_001110001110: DATA = 12'b000000100000;
            14'b10_001110001111: DATA = 12'b000000011111;
            14'b10_001110010000: DATA = 12'b000000011111;
            14'b10_001110010001: DATA = 12'b000000011110;
            14'b10_001110010010: DATA = 12'b000000011110;
            14'b10_001110010011: DATA = 12'b000000011101;
            14'b10_001110010100: DATA = 12'b000000011101;
            14'b10_001110010101: DATA = 12'b000000011100;
            14'b10_001110010110: DATA = 12'b000000011100;
            14'b10_001110010111: DATA = 12'b000000011011;
            14'b10_001110011000: DATA = 12'b000000011010;
            14'b10_001110011001: DATA = 12'b000000011010;
            14'b10_001110011010: DATA = 12'b000000011010;
            14'b10_001110011011: DATA = 12'b000000011001;
            14'b10_001110011100: DATA = 12'b000000011001;
            14'b10_001110011101: DATA = 12'b000000011000;
            14'b10_001110011110: DATA = 12'b000000011000;
            14'b10_001110011111: DATA = 12'b000000010111;
            14'b10_001110100000: DATA = 12'b000000010111;
            14'b10_001110100001: DATA = 12'b000000010110;
            14'b10_001110100010: DATA = 12'b000000010110;
            14'b10_001110100011: DATA = 12'b000000010101;
            14'b10_001110100100: DATA = 12'b000000010101;
            14'b10_001110100101: DATA = 12'b000000010100;
            14'b10_001110100110: DATA = 12'b000000010100;
            14'b10_001110100111: DATA = 12'b000000010100;
            14'b10_001110101000: DATA = 12'b000000010011;
            14'b10_001110101001: DATA = 12'b000000010011;
            14'b10_001110101010: DATA = 12'b000000010010;
            14'b10_001110101011: DATA = 12'b000000010010;
            14'b10_001110101100: DATA = 12'b000000010001;
            14'b10_001110101101: DATA = 12'b000000010001;
            14'b10_001110101110: DATA = 12'b000000010001;
            14'b10_001110101111: DATA = 12'b000000010000;
            14'b10_001110110000: DATA = 12'b000000010000;
            14'b10_001110110001: DATA = 12'b000000010000;
            14'b10_001110110010: DATA = 12'b000000001111;
            14'b10_001110110011: DATA = 12'b000000001111;
            14'b10_001110110100: DATA = 12'b000000001110;
            14'b10_001110110101: DATA = 12'b000000001110;
            14'b10_001110110110: DATA = 12'b000000001110;
            14'b10_001110110111: DATA = 12'b000000001101;
            14'b10_001110111000: DATA = 12'b000000001101;
            14'b10_001110111001: DATA = 12'b000000001101;
            14'b10_001110111010: DATA = 12'b000000001100;
            14'b10_001110111011: DATA = 12'b000000001100;
            14'b10_001110111100: DATA = 12'b000000001100;
            14'b10_001110111101: DATA = 12'b000000001011;
            14'b10_001110111110: DATA = 12'b000000001011;
            14'b10_001110111111: DATA = 12'b000000001011;
            14'b10_001111000000: DATA = 12'b000000001010;
            14'b10_001111000001: DATA = 12'b000000001010;
            14'b10_001111000010: DATA = 12'b000000001010;
            14'b10_001111000011: DATA = 12'b000000001001;
            14'b10_001111000100: DATA = 12'b000000001001;
            14'b10_001111000101: DATA = 12'b000000001001;
            14'b10_001111000110: DATA = 12'b000000001001;
            14'b10_001111000111: DATA = 12'b000000001000;
            14'b10_001111001000: DATA = 12'b000000001000;
            14'b10_001111001001: DATA = 12'b000000001000;
            14'b10_001111001010: DATA = 12'b000000001000;
            14'b10_001111001011: DATA = 12'b000000000111;
            14'b10_001111001100: DATA = 12'b000000000111;
            14'b10_001111001101: DATA = 12'b000000000111;
            14'b10_001111001110: DATA = 12'b000000000111;
            14'b10_001111001111: DATA = 12'b000000000110;
            14'b10_001111010000: DATA = 12'b000000000110;
            14'b10_001111010001: DATA = 12'b000000000110;
            14'b10_001111010010: DATA = 12'b000000000110;
            14'b10_001111010011: DATA = 12'b000000000101;
            14'b10_001111010100: DATA = 12'b000000000101;
            14'b10_001111010101: DATA = 12'b000000000101;
            14'b10_001111010110: DATA = 12'b000000000101;
            14'b10_001111010111: DATA = 12'b000000000101;
            14'b10_001111011000: DATA = 12'b000000000100;
            14'b10_001111011001: DATA = 12'b000000000100;
            14'b10_001111011010: DATA = 12'b000000000100;
            14'b10_001111011011: DATA = 12'b000000000100;
            14'b10_001111011100: DATA = 12'b000000000100;
            14'b10_001111011101: DATA = 12'b000000000011;
            14'b10_001111011110: DATA = 12'b000000000011;
            14'b10_001111011111: DATA = 12'b000000000011;
            14'b10_001111100000: DATA = 12'b000000000011;
            14'b10_001111100001: DATA = 12'b000000000011;
            14'b10_001111100010: DATA = 12'b000000000011;
            14'b10_001111100011: DATA = 12'b000000000011;
            14'b10_001111100100: DATA = 12'b000000000010;
            14'b10_001111100101: DATA = 12'b000000000010;
            14'b10_001111100110: DATA = 12'b000000000010;
            14'b10_001111100111: DATA = 12'b000000000010;
            14'b10_001111101000: DATA = 12'b000000000010;
            14'b10_001111101001: DATA = 12'b000000000010;
            14'b10_001111101010: DATA = 12'b000000000010;
            14'b10_001111101011: DATA = 12'b000000000010;
            14'b10_001111101100: DATA = 12'b000000000001;
            14'b10_001111101101: DATA = 12'b000000000001;
            14'b10_001111101110: DATA = 12'b000000000001;
            14'b10_001111101111: DATA = 12'b000000000001;
            14'b10_001111110000: DATA = 12'b000000000001;
            14'b10_001111110001: DATA = 12'b000000000001;
            14'b10_001111110010: DATA = 12'b000000000001;
            14'b10_001111110011: DATA = 12'b000000000001;
            14'b10_001111110100: DATA = 12'b000000000001;
            14'b10_001111110101: DATA = 12'b000000000001;
            14'b10_001111110110: DATA = 12'b000000000001;
            14'b10_001111110111: DATA = 12'b000000000001;
            14'b10_001111111000: DATA = 12'b000000000001;
            14'b10_001111111001: DATA = 12'b000000000001;
            14'b10_001111111010: DATA = 12'b000000000001;
            14'b10_001111111011: DATA = 12'b000000000001;
            14'b10_001111111100: DATA = 12'b000000000001;
            14'b10_001111111101: DATA = 12'b000000000001;
            14'b10_001111111110: DATA = 12'b000000000001;
            14'b10_001111111111: DATA = 12'b000000000001;
            14'b10_010000000000: DATA = 12'b000000000001;
            14'b10_010000000001: DATA = 12'b000000000001;
            14'b10_010000000010: DATA = 12'b000000000001;
            14'b10_010000000011: DATA = 12'b000000000001;
            14'b10_010000000100: DATA = 12'b000000000001;
            14'b10_010000000101: DATA = 12'b000000000001;
            14'b10_010000000110: DATA = 12'b000000000001;
            14'b10_010000000111: DATA = 12'b000000000001;
            14'b10_010000001000: DATA = 12'b000000000001;
            14'b10_010000001001: DATA = 12'b000000000001;
            14'b10_010000001010: DATA = 12'b000000000001;
            14'b10_010000001011: DATA = 12'b000000000001;
            14'b10_010000001100: DATA = 12'b000000000001;
            14'b10_010000001101: DATA = 12'b000000000001;
            14'b10_010000001110: DATA = 12'b000000000001;
            14'b10_010000001111: DATA = 12'b000000000001;
            14'b10_010000010000: DATA = 12'b000000000001;
            14'b10_010000010001: DATA = 12'b000000000001;
            14'b10_010000010010: DATA = 12'b000000000001;
            14'b10_010000010011: DATA = 12'b000000000001;
            14'b10_010000010100: DATA = 12'b000000000001;
            14'b10_010000010101: DATA = 12'b000000000010;
            14'b10_010000010110: DATA = 12'b000000000010;
            14'b10_010000010111: DATA = 12'b000000000010;
            14'b10_010000011000: DATA = 12'b000000000010;
            14'b10_010000011001: DATA = 12'b000000000010;
            14'b10_010000011010: DATA = 12'b000000000010;
            14'b10_010000011011: DATA = 12'b000000000010;
            14'b10_010000011100: DATA = 12'b000000000010;
            14'b10_010000011101: DATA = 12'b000000000011;
            14'b10_010000011110: DATA = 12'b000000000011;
            14'b10_010000011111: DATA = 12'b000000000011;
            14'b10_010000100000: DATA = 12'b000000000011;
            14'b10_010000100001: DATA = 12'b000000000011;
            14'b10_010000100010: DATA = 12'b000000000011;
            14'b10_010000100011: DATA = 12'b000000000011;
            14'b10_010000100100: DATA = 12'b000000000100;
            14'b10_010000100101: DATA = 12'b000000000100;
            14'b10_010000100110: DATA = 12'b000000000100;
            14'b10_010000100111: DATA = 12'b000000000100;
            14'b10_010000101000: DATA = 12'b000000000100;
            14'b10_010000101001: DATA = 12'b000000000101;
            14'b10_010000101010: DATA = 12'b000000000101;
            14'b10_010000101011: DATA = 12'b000000000101;
            14'b10_010000101100: DATA = 12'b000000000101;
            14'b10_010000101101: DATA = 12'b000000000101;
            14'b10_010000101110: DATA = 12'b000000000110;
            14'b10_010000101111: DATA = 12'b000000000110;
            14'b10_010000110000: DATA = 12'b000000000110;
            14'b10_010000110001: DATA = 12'b000000000110;
            14'b10_010000110010: DATA = 12'b000000000111;
            14'b10_010000110011: DATA = 12'b000000000111;
            14'b10_010000110100: DATA = 12'b000000000111;
            14'b10_010000110101: DATA = 12'b000000000111;
            14'b10_010000110110: DATA = 12'b000000001000;
            14'b10_010000110111: DATA = 12'b000000001000;
            14'b10_010000111000: DATA = 12'b000000001000;
            14'b10_010000111001: DATA = 12'b000000001000;
            14'b10_010000111010: DATA = 12'b000000001001;
            14'b10_010000111011: DATA = 12'b000000001001;
            14'b10_010000111100: DATA = 12'b000000001001;
            14'b10_010000111101: DATA = 12'b000000001001;
            14'b10_010000111110: DATA = 12'b000000001010;
            14'b10_010000111111: DATA = 12'b000000001010;
            14'b10_010001000000: DATA = 12'b000000001010;
            14'b10_010001000001: DATA = 12'b000000001011;
            14'b10_010001000010: DATA = 12'b000000001011;
            14'b10_010001000011: DATA = 12'b000000001011;
            14'b10_010001000100: DATA = 12'b000000001100;
            14'b10_010001000101: DATA = 12'b000000001100;
            14'b10_010001000110: DATA = 12'b000000001100;
            14'b10_010001000111: DATA = 12'b000000001101;
            14'b10_010001001000: DATA = 12'b000000001101;
            14'b10_010001001001: DATA = 12'b000000001101;
            14'b10_010001001010: DATA = 12'b000000001110;
            14'b10_010001001011: DATA = 12'b000000001110;
            14'b10_010001001100: DATA = 12'b000000001110;
            14'b10_010001001101: DATA = 12'b000000001111;
            14'b10_010001001110: DATA = 12'b000000001111;
            14'b10_010001001111: DATA = 12'b000000010000;
            14'b10_010001010000: DATA = 12'b000000010000;
            14'b10_010001010001: DATA = 12'b000000010000;
            14'b10_010001010010: DATA = 12'b000000010001;
            14'b10_010001010011: DATA = 12'b000000010001;
            14'b10_010001010100: DATA = 12'b000000010001;
            14'b10_010001010101: DATA = 12'b000000010010;
            14'b10_010001010110: DATA = 12'b000000010010;
            14'b10_010001010111: DATA = 12'b000000010011;
            14'b10_010001011000: DATA = 12'b000000010011;
            14'b10_010001011001: DATA = 12'b000000010100;
            14'b10_010001011010: DATA = 12'b000000010100;
            14'b10_010001011011: DATA = 12'b000000010100;
            14'b10_010001011100: DATA = 12'b000000010101;
            14'b10_010001011101: DATA = 12'b000000010101;
            14'b10_010001011110: DATA = 12'b000000010110;
            14'b10_010001011111: DATA = 12'b000000010110;
            14'b10_010001100000: DATA = 12'b000000010111;
            14'b10_010001100001: DATA = 12'b000000010111;
            14'b10_010001100010: DATA = 12'b000000011000;
            14'b10_010001100011: DATA = 12'b000000011000;
            14'b10_010001100100: DATA = 12'b000000011001;
            14'b10_010001100101: DATA = 12'b000000011001;
            14'b10_010001100110: DATA = 12'b000000011010;
            14'b10_010001100111: DATA = 12'b000000011010;
            14'b10_010001101000: DATA = 12'b000000011010;
            14'b10_010001101001: DATA = 12'b000000011011;
            14'b10_010001101010: DATA = 12'b000000011100;
            14'b10_010001101011: DATA = 12'b000000011100;
            14'b10_010001101100: DATA = 12'b000000011101;
            14'b10_010001101101: DATA = 12'b000000011101;
            14'b10_010001101110: DATA = 12'b000000011110;
            14'b10_010001101111: DATA = 12'b000000011110;
            14'b10_010001110000: DATA = 12'b000000011111;
            14'b10_010001110001: DATA = 12'b000000011111;
            14'b10_010001110010: DATA = 12'b000000100000;
            14'b10_010001110011: DATA = 12'b000000100000;
            14'b10_010001110100: DATA = 12'b000000100001;
            14'b10_010001110101: DATA = 12'b000000100001;
            14'b10_010001110110: DATA = 12'b000000100010;
            14'b10_010001110111: DATA = 12'b000000100011;
            14'b10_010001111000: DATA = 12'b000000100011;
            14'b10_010001111001: DATA = 12'b000000100100;
            14'b10_010001111010: DATA = 12'b000000100100;
            14'b10_010001111011: DATA = 12'b000000100101;
            14'b10_010001111100: DATA = 12'b000000100101;
            14'b10_010001111101: DATA = 12'b000000100110;
            14'b10_010001111110: DATA = 12'b000000100111;
            14'b10_010001111111: DATA = 12'b000000100111;
            14'b10_010010000000: DATA = 12'b000000101000;
            14'b10_010010000001: DATA = 12'b000000101000;
            14'b10_010010000010: DATA = 12'b000000101001;
            14'b10_010010000011: DATA = 12'b000000101010;
            14'b10_010010000100: DATA = 12'b000000101010;
            14'b10_010010000101: DATA = 12'b000000101011;
            14'b10_010010000110: DATA = 12'b000000101100;
            14'b10_010010000111: DATA = 12'b000000101100;
            14'b10_010010001000: DATA = 12'b000000101101;
            14'b10_010010001001: DATA = 12'b000000101110;
            14'b10_010010001010: DATA = 12'b000000101110;
            14'b10_010010001011: DATA = 12'b000000101111;
            14'b10_010010001100: DATA = 12'b000000110000;
            14'b10_010010001101: DATA = 12'b000000110000;
            14'b10_010010001110: DATA = 12'b000000110001;
            14'b10_010010001111: DATA = 12'b000000110010;
            14'b10_010010010000: DATA = 12'b000000110010;
            14'b10_010010010001: DATA = 12'b000000110011;
            14'b10_010010010010: DATA = 12'b000000110100;
            14'b10_010010010011: DATA = 12'b000000110100;
            14'b10_010010010100: DATA = 12'b000000110101;
            14'b10_010010010101: DATA = 12'b000000110110;
            14'b10_010010010110: DATA = 12'b000000110110;
            14'b10_010010010111: DATA = 12'b000000110111;
            14'b10_010010011000: DATA = 12'b000000111000;
            14'b10_010010011001: DATA = 12'b000000111001;
            14'b10_010010011010: DATA = 12'b000000111001;
            14'b10_010010011011: DATA = 12'b000000111010;
            14'b10_010010011100: DATA = 12'b000000111011;
            14'b10_010010011101: DATA = 12'b000000111100;
            14'b10_010010011110: DATA = 12'b000000111100;
            14'b10_010010011111: DATA = 12'b000000111101;
            14'b10_010010100000: DATA = 12'b000000111110;
            14'b10_010010100001: DATA = 12'b000000111111;
            14'b10_010010100010: DATA = 12'b000000111111;
            14'b10_010010100011: DATA = 12'b000001000000;
            14'b10_010010100100: DATA = 12'b000001000001;
            14'b10_010010100101: DATA = 12'b000001000010;
            14'b10_010010100110: DATA = 12'b000001000011;
            14'b10_010010100111: DATA = 12'b000001000011;
            14'b10_010010101000: DATA = 12'b000001000100;
            14'b10_010010101001: DATA = 12'b000001000101;
            14'b10_010010101010: DATA = 12'b000001000110;
            14'b10_010010101011: DATA = 12'b000001000111;
            14'b10_010010101100: DATA = 12'b000001000111;
            14'b10_010010101101: DATA = 12'b000001001000;
            14'b10_010010101110: DATA = 12'b000001001001;
            14'b10_010010101111: DATA = 12'b000001001010;
            14'b10_010010110000: DATA = 12'b000001001011;
            14'b10_010010110001: DATA = 12'b000001001011;
            14'b10_010010110010: DATA = 12'b000001001100;
            14'b10_010010110011: DATA = 12'b000001001101;
            14'b10_010010110100: DATA = 12'b000001001110;
            14'b10_010010110101: DATA = 12'b000001001111;
            14'b10_010010110110: DATA = 12'b000001010000;
            14'b10_010010110111: DATA = 12'b000001010001;
            14'b10_010010111000: DATA = 12'b000001010001;
            14'b10_010010111001: DATA = 12'b000001010010;
            14'b10_010010111010: DATA = 12'b000001010011;
            14'b10_010010111011: DATA = 12'b000001010100;
            14'b10_010010111100: DATA = 12'b000001010101;
            14'b10_010010111101: DATA = 12'b000001010110;
            14'b10_010010111110: DATA = 12'b000001010111;
            14'b10_010010111111: DATA = 12'b000001011000;
            14'b10_010011000000: DATA = 12'b000001011001;
            14'b10_010011000001: DATA = 12'b000001011010;
            14'b10_010011000010: DATA = 12'b000001011010;
            14'b10_010011000011: DATA = 12'b000001011011;
            14'b10_010011000100: DATA = 12'b000001011100;
            14'b10_010011000101: DATA = 12'b000001011101;
            14'b10_010011000110: DATA = 12'b000001011110;
            14'b10_010011000111: DATA = 12'b000001011111;
            14'b10_010011001000: DATA = 12'b000001100000;
            14'b10_010011001001: DATA = 12'b000001100001;
            14'b10_010011001010: DATA = 12'b000001100010;
            14'b10_010011001011: DATA = 12'b000001100011;
            14'b10_010011001100: DATA = 12'b000001100100;
            14'b10_010011001101: DATA = 12'b000001100101;
            14'b10_010011001110: DATA = 12'b000001100110;
            14'b10_010011001111: DATA = 12'b000001100111;
            14'b10_010011010000: DATA = 12'b000001101000;
            14'b10_010011010001: DATA = 12'b000001101001;
            14'b10_010011010010: DATA = 12'b000001101010;
            14'b10_010011010011: DATA = 12'b000001101011;
            14'b10_010011010100: DATA = 12'b000001101100;
            14'b10_010011010101: DATA = 12'b000001101101;
            14'b10_010011010110: DATA = 12'b000001101110;
            14'b10_010011010111: DATA = 12'b000001101111;
            14'b10_010011011000: DATA = 12'b000001110000;
            14'b10_010011011001: DATA = 12'b000001110001;
            14'b10_010011011010: DATA = 12'b000001110010;
            14'b10_010011011011: DATA = 12'b000001110011;
            14'b10_010011011100: DATA = 12'b000001110100;
            14'b10_010011011101: DATA = 12'b000001110101;
            14'b10_010011011110: DATA = 12'b000001110110;
            14'b10_010011011111: DATA = 12'b000001110111;
            14'b10_010011100000: DATA = 12'b000001111000;
            14'b10_010011100001: DATA = 12'b000001111001;
            14'b10_010011100010: DATA = 12'b000001111010;
            14'b10_010011100011: DATA = 12'b000001111011;
            14'b10_010011100100: DATA = 12'b000001111100;
            14'b10_010011100101: DATA = 12'b000001111110;
            14'b10_010011100110: DATA = 12'b000001111111;
            14'b10_010011100111: DATA = 12'b000010000000;
            14'b10_010011101000: DATA = 12'b000010000001;
            14'b10_010011101001: DATA = 12'b000010000010;
            14'b10_010011101010: DATA = 12'b000010000011;
            14'b10_010011101011: DATA = 12'b000010000100;
            14'b10_010011101100: DATA = 12'b000010000101;
            14'b10_010011101101: DATA = 12'b000010000110;
            14'b10_010011101110: DATA = 12'b000010000111;
            14'b10_010011101111: DATA = 12'b000010001001;
            14'b10_010011110000: DATA = 12'b000010001010;
            14'b10_010011110001: DATA = 12'b000010001011;
            14'b10_010011110010: DATA = 12'b000010001100;
            14'b10_010011110011: DATA = 12'b000010001101;
            14'b10_010011110100: DATA = 12'b000010001110;
            14'b10_010011110101: DATA = 12'b000010001111;
            14'b10_010011110110: DATA = 12'b000010010001;
            14'b10_010011110111: DATA = 12'b000010010010;
            14'b10_010011111000: DATA = 12'b000010010011;
            14'b10_010011111001: DATA = 12'b000010010100;
            14'b10_010011111010: DATA = 12'b000010010101;
            14'b10_010011111011: DATA = 12'b000010010110;
            14'b10_010011111100: DATA = 12'b000010011000;
            14'b10_010011111101: DATA = 12'b000010011001;
            14'b10_010011111110: DATA = 12'b000010011010;
            14'b10_010011111111: DATA = 12'b000010011011;
            14'b10_010100000000: DATA = 12'b000010011100;
            14'b10_010100000001: DATA = 12'b000010011110;
            14'b10_010100000010: DATA = 12'b000010011111;
            14'b10_010100000011: DATA = 12'b000010100000;
            14'b10_010100000100: DATA = 12'b000010100001;
            14'b10_010100000101: DATA = 12'b000010100010;
            14'b10_010100000110: DATA = 12'b000010100100;
            14'b10_010100000111: DATA = 12'b000010100101;
            14'b10_010100001000: DATA = 12'b000010100110;
            14'b10_010100001001: DATA = 12'b000010100111;
            14'b10_010100001010: DATA = 12'b000010101001;
            14'b10_010100001011: DATA = 12'b000010101010;
            14'b10_010100001100: DATA = 12'b000010101011;
            14'b10_010100001101: DATA = 12'b000010101100;
            14'b10_010100001110: DATA = 12'b000010101110;
            14'b10_010100001111: DATA = 12'b000010101111;
            14'b10_010100010000: DATA = 12'b000010110000;
            14'b10_010100010001: DATA = 12'b000010110001;
            14'b10_010100010010: DATA = 12'b000010110011;
            14'b10_010100010011: DATA = 12'b000010110100;
            14'b10_010100010100: DATA = 12'b000010110101;
            14'b10_010100010101: DATA = 12'b000010110111;
            14'b10_010100010110: DATA = 12'b000010111000;
            14'b10_010100010111: DATA = 12'b000010111001;
            14'b10_010100011000: DATA = 12'b000010111010;
            14'b10_010100011001: DATA = 12'b000010111100;
            14'b10_010100011010: DATA = 12'b000010111101;
            14'b10_010100011011: DATA = 12'b000010111110;
            14'b10_010100011100: DATA = 12'b000011000000;
            14'b10_010100011101: DATA = 12'b000011000001;
            14'b10_010100011110: DATA = 12'b000011000010;
            14'b10_010100011111: DATA = 12'b000011000100;
            14'b10_010100100000: DATA = 12'b000011000101;
            14'b10_010100100001: DATA = 12'b000011000110;
            14'b10_010100100010: DATA = 12'b000011001000;
            14'b10_010100100011: DATA = 12'b000011001001;
            14'b10_010100100100: DATA = 12'b000011001010;
            14'b10_010100100101: DATA = 12'b000011001100;
            14'b10_010100100110: DATA = 12'b000011001101;
            14'b10_010100100111: DATA = 12'b000011001111;
            14'b10_010100101000: DATA = 12'b000011010000;
            14'b10_010100101001: DATA = 12'b000011010001;
            14'b10_010100101010: DATA = 12'b000011010011;
            14'b10_010100101011: DATA = 12'b000011010100;
            14'b10_010100101100: DATA = 12'b000011010101;
            14'b10_010100101101: DATA = 12'b000011010111;
            14'b10_010100101110: DATA = 12'b000011011000;
            14'b10_010100101111: DATA = 12'b000011011010;
            14'b10_010100110000: DATA = 12'b000011011011;
            14'b10_010100110001: DATA = 12'b000011011100;
            14'b10_010100110010: DATA = 12'b000011011110;
            14'b10_010100110011: DATA = 12'b000011011111;
            14'b10_010100110100: DATA = 12'b000011100001;
            14'b10_010100110101: DATA = 12'b000011100010;
            14'b10_010100110110: DATA = 12'b000011100100;
            14'b10_010100110111: DATA = 12'b000011100101;
            14'b10_010100111000: DATA = 12'b000011100111;
            14'b10_010100111001: DATA = 12'b000011101000;
            14'b10_010100111010: DATA = 12'b000011101001;
            14'b10_010100111011: DATA = 12'b000011101011;
            14'b10_010100111100: DATA = 12'b000011101100;
            14'b10_010100111101: DATA = 12'b000011101110;
            14'b10_010100111110: DATA = 12'b000011101111;
            14'b10_010100111111: DATA = 12'b000011110001;
            14'b10_010101000000: DATA = 12'b000011110010;
            14'b10_010101000001: DATA = 12'b000011110100;
            14'b10_010101000010: DATA = 12'b000011110101;
            14'b10_010101000011: DATA = 12'b000011110111;
            14'b10_010101000100: DATA = 12'b000011111000;
            14'b10_010101000101: DATA = 12'b000011111010;
            14'b10_010101000110: DATA = 12'b000011111011;
            14'b10_010101000111: DATA = 12'b000011111101;
            14'b10_010101001000: DATA = 12'b000011111110;
            14'b10_010101001001: DATA = 12'b000100000000;
            14'b10_010101001010: DATA = 12'b000100000001;
            14'b10_010101001011: DATA = 12'b000100000011;
            14'b10_010101001100: DATA = 12'b000100000100;
            14'b10_010101001101: DATA = 12'b000100000110;
            14'b10_010101001110: DATA = 12'b000100000111;
            14'b10_010101001111: DATA = 12'b000100001001;
            14'b10_010101010000: DATA = 12'b000100001010;
            14'b10_010101010001: DATA = 12'b000100001100;
            14'b10_010101010010: DATA = 12'b000100001110;
            14'b10_010101010011: DATA = 12'b000100001111;
            14'b10_010101010100: DATA = 12'b000100010001;
            14'b10_010101010101: DATA = 12'b000100010010;
            14'b10_010101010110: DATA = 12'b000100010100;
            14'b10_010101010111: DATA = 12'b000100010101;
            14'b10_010101011000: DATA = 12'b000100010111;
            14'b10_010101011001: DATA = 12'b000100011001;
            14'b10_010101011010: DATA = 12'b000100011010;
            14'b10_010101011011: DATA = 12'b000100011100;
            14'b10_010101011100: DATA = 12'b000100011101;
            14'b10_010101011101: DATA = 12'b000100011111;
            14'b10_010101011110: DATA = 12'b000100100001;
            14'b10_010101011111: DATA = 12'b000100100010;
            14'b10_010101100000: DATA = 12'b000100100100;
            14'b10_010101100001: DATA = 12'b000100100101;
            14'b10_010101100010: DATA = 12'b000100100111;
            14'b10_010101100011: DATA = 12'b000100101001;
            14'b10_010101100100: DATA = 12'b000100101010;
            14'b10_010101100101: DATA = 12'b000100101100;
            14'b10_010101100110: DATA = 12'b000100101101;
            14'b10_010101100111: DATA = 12'b000100101111;
            14'b10_010101101000: DATA = 12'b000100110001;
            14'b10_010101101001: DATA = 12'b000100110010;
            14'b10_010101101010: DATA = 12'b000100110100;
            14'b10_010101101011: DATA = 12'b000100110110;
            14'b10_010101101100: DATA = 12'b000100110111;
            14'b10_010101101101: DATA = 12'b000100111001;
            14'b10_010101101110: DATA = 12'b000100111011;
            14'b10_010101101111: DATA = 12'b000100111100;
            14'b10_010101110000: DATA = 12'b000100111110;
            14'b10_010101110001: DATA = 12'b000101000000;
            14'b10_010101110010: DATA = 12'b000101000001;
            14'b10_010101110011: DATA = 12'b000101000011;
            14'b10_010101110100: DATA = 12'b000101000101;
            14'b10_010101110101: DATA = 12'b000101000111;
            14'b10_010101110110: DATA = 12'b000101001000;
            14'b10_010101110111: DATA = 12'b000101001010;
            14'b10_010101111000: DATA = 12'b000101001100;
            14'b10_010101111001: DATA = 12'b000101001101;
            14'b10_010101111010: DATA = 12'b000101001111;
            14'b10_010101111011: DATA = 12'b000101010001;
            14'b10_010101111100: DATA = 12'b000101010011;
            14'b10_010101111101: DATA = 12'b000101010100;
            14'b10_010101111110: DATA = 12'b000101010110;
            14'b10_010101111111: DATA = 12'b000101011000;
            14'b10_010110000000: DATA = 12'b000101011001;
            14'b10_010110000001: DATA = 12'b000101011011;
            14'b10_010110000010: DATA = 12'b000101011101;
            14'b10_010110000011: DATA = 12'b000101011111;
            14'b10_010110000100: DATA = 12'b000101100000;
            14'b10_010110000101: DATA = 12'b000101100010;
            14'b10_010110000110: DATA = 12'b000101100100;
            14'b10_010110000111: DATA = 12'b000101100110;
            14'b10_010110001000: DATA = 12'b000101101000;
            14'b10_010110001001: DATA = 12'b000101101001;
            14'b10_010110001010: DATA = 12'b000101101011;
            14'b10_010110001011: DATA = 12'b000101101101;
            14'b10_010110001100: DATA = 12'b000101101111;
            14'b10_010110001101: DATA = 12'b000101110000;
            14'b10_010110001110: DATA = 12'b000101110010;
            14'b10_010110001111: DATA = 12'b000101110100;
            14'b10_010110010000: DATA = 12'b000101110110;
            14'b10_010110010001: DATA = 12'b000101111000;
            14'b10_010110010010: DATA = 12'b000101111010;
            14'b10_010110010011: DATA = 12'b000101111011;
            14'b10_010110010100: DATA = 12'b000101111101;
            14'b10_010110010101: DATA = 12'b000101111111;
            14'b10_010110010110: DATA = 12'b000110000001;
            14'b10_010110010111: DATA = 12'b000110000011;
            14'b10_010110011000: DATA = 12'b000110000100;
            14'b10_010110011001: DATA = 12'b000110000110;
            14'b10_010110011010: DATA = 12'b000110001000;
            14'b10_010110011011: DATA = 12'b000110001010;
            14'b10_010110011100: DATA = 12'b000110001100;
            14'b10_010110011101: DATA = 12'b000110001110;
            14'b10_010110011110: DATA = 12'b000110010000;
            14'b10_010110011111: DATA = 12'b000110010001;
            14'b10_010110100000: DATA = 12'b000110010011;
            14'b10_010110100001: DATA = 12'b000110010101;
            14'b10_010110100010: DATA = 12'b000110010111;
            14'b10_010110100011: DATA = 12'b000110011001;
            14'b10_010110100100: DATA = 12'b000110011011;
            14'b10_010110100101: DATA = 12'b000110011101;
            14'b10_010110100110: DATA = 12'b000110011111;
            14'b10_010110100111: DATA = 12'b000110100001;
            14'b10_010110101000: DATA = 12'b000110100010;
            14'b10_010110101001: DATA = 12'b000110100100;
            14'b10_010110101010: DATA = 12'b000110100110;
            14'b10_010110101011: DATA = 12'b000110101000;
            14'b10_010110101100: DATA = 12'b000110101010;
            14'b10_010110101101: DATA = 12'b000110101100;
            14'b10_010110101110: DATA = 12'b000110101110;
            14'b10_010110101111: DATA = 12'b000110110000;
            14'b10_010110110000: DATA = 12'b000110110010;
            14'b10_010110110001: DATA = 12'b000110110100;
            14'b10_010110110010: DATA = 12'b000110110110;
            14'b10_010110110011: DATA = 12'b000110111000;
            14'b10_010110110100: DATA = 12'b000110111010;
            14'b10_010110110101: DATA = 12'b000110111011;
            14'b10_010110110110: DATA = 12'b000110111101;
            14'b10_010110110111: DATA = 12'b000110111111;
            14'b10_010110111000: DATA = 12'b000111000001;
            14'b10_010110111001: DATA = 12'b000111000011;
            14'b10_010110111010: DATA = 12'b000111000101;
            14'b10_010110111011: DATA = 12'b000111000111;
            14'b10_010110111100: DATA = 12'b000111001001;
            14'b10_010110111101: DATA = 12'b000111001011;
            14'b10_010110111110: DATA = 12'b000111001101;
            14'b10_010110111111: DATA = 12'b000111001111;
            14'b10_010111000000: DATA = 12'b000111010001;
            14'b10_010111000001: DATA = 12'b000111010011;
            14'b10_010111000010: DATA = 12'b000111010101;
            14'b10_010111000011: DATA = 12'b000111010111;
            14'b10_010111000100: DATA = 12'b000111011001;
            14'b10_010111000101: DATA = 12'b000111011011;
            14'b10_010111000110: DATA = 12'b000111011101;
            14'b10_010111000111: DATA = 12'b000111011111;
            14'b10_010111001000: DATA = 12'b000111100001;
            14'b10_010111001001: DATA = 12'b000111100011;
            14'b10_010111001010: DATA = 12'b000111100101;
            14'b10_010111001011: DATA = 12'b000111100111;
            14'b10_010111001100: DATA = 12'b000111101001;
            14'b10_010111001101: DATA = 12'b000111101011;
            14'b10_010111001110: DATA = 12'b000111101101;
            14'b10_010111001111: DATA = 12'b000111101111;
            14'b10_010111010000: DATA = 12'b000111110001;
            14'b10_010111010001: DATA = 12'b000111110100;
            14'b10_010111010010: DATA = 12'b000111110110;
            14'b10_010111010011: DATA = 12'b000111111000;
            14'b10_010111010100: DATA = 12'b000111111010;
            14'b10_010111010101: DATA = 12'b000111111100;
            14'b10_010111010110: DATA = 12'b000111111110;
            14'b10_010111010111: DATA = 12'b001000000000;
            14'b10_010111011000: DATA = 12'b001000000010;
            14'b10_010111011001: DATA = 12'b001000000100;
            14'b10_010111011010: DATA = 12'b001000000110;
            14'b10_010111011011: DATA = 12'b001000001000;
            14'b10_010111011100: DATA = 12'b001000001010;
            14'b10_010111011101: DATA = 12'b001000001100;
            14'b10_010111011110: DATA = 12'b001000001111;
            14'b10_010111011111: DATA = 12'b001000010001;
            14'b10_010111100000: DATA = 12'b001000010011;
            14'b10_010111100001: DATA = 12'b001000010101;
            14'b10_010111100010: DATA = 12'b001000010111;
            14'b10_010111100011: DATA = 12'b001000011001;
            14'b10_010111100100: DATA = 12'b001000011011;
            14'b10_010111100101: DATA = 12'b001000011101;
            14'b10_010111100110: DATA = 12'b001000011111;
            14'b10_010111100111: DATA = 12'b001000100010;
            14'b10_010111101000: DATA = 12'b001000100100;
            14'b10_010111101001: DATA = 12'b001000100110;
            14'b10_010111101010: DATA = 12'b001000101000;
            14'b10_010111101011: DATA = 12'b001000101010;
            14'b10_010111101100: DATA = 12'b001000101100;
            14'b10_010111101101: DATA = 12'b001000101110;
            14'b10_010111101110: DATA = 12'b001000110001;
            14'b10_010111101111: DATA = 12'b001000110011;
            14'b10_010111110000: DATA = 12'b001000110101;
            14'b10_010111110001: DATA = 12'b001000110111;
            14'b10_010111110010: DATA = 12'b001000111001;
            14'b10_010111110011: DATA = 12'b001000111011;
            14'b10_010111110100: DATA = 12'b001000111110;
            14'b10_010111110101: DATA = 12'b001001000000;
            14'b10_010111110110: DATA = 12'b001001000010;
            14'b10_010111110111: DATA = 12'b001001000100;
            14'b10_010111111000: DATA = 12'b001001000110;
            14'b10_010111111001: DATA = 12'b001001001001;
            14'b10_010111111010: DATA = 12'b001001001011;
            14'b10_010111111011: DATA = 12'b001001001101;
            14'b10_010111111100: DATA = 12'b001001001111;
            14'b10_010111111101: DATA = 12'b001001010001;
            14'b10_010111111110: DATA = 12'b001001010100;
            14'b10_010111111111: DATA = 12'b001001010110;
            14'b10_011000000000: DATA = 12'b001001011000;
            14'b10_011000000001: DATA = 12'b001001011010;
            14'b10_011000000010: DATA = 12'b001001011100;
            14'b10_011000000011: DATA = 12'b001001011111;
            14'b10_011000000100: DATA = 12'b001001100001;
            14'b10_011000000101: DATA = 12'b001001100011;
            14'b10_011000000110: DATA = 12'b001001100101;
            14'b10_011000000111: DATA = 12'b001001101000;
            14'b10_011000001000: DATA = 12'b001001101010;
            14'b10_011000001001: DATA = 12'b001001101100;
            14'b10_011000001010: DATA = 12'b001001101110;
            14'b10_011000001011: DATA = 12'b001001110001;
            14'b10_011000001100: DATA = 12'b001001110011;
            14'b10_011000001101: DATA = 12'b001001110101;
            14'b10_011000001110: DATA = 12'b001001110111;
            14'b10_011000001111: DATA = 12'b001001111010;
            14'b10_011000010000: DATA = 12'b001001111100;
            14'b10_011000010001: DATA = 12'b001001111110;
            14'b10_011000010010: DATA = 12'b001010000001;
            14'b10_011000010011: DATA = 12'b001010000011;
            14'b10_011000010100: DATA = 12'b001010000101;
            14'b10_011000010101: DATA = 12'b001010000111;
            14'b10_011000010110: DATA = 12'b001010001010;
            14'b10_011000010111: DATA = 12'b001010001100;
            14'b10_011000011000: DATA = 12'b001010001110;
            14'b10_011000011001: DATA = 12'b001010010001;
            14'b10_011000011010: DATA = 12'b001010010011;
            14'b10_011000011011: DATA = 12'b001010010101;
            14'b10_011000011100: DATA = 12'b001010011000;
            14'b10_011000011101: DATA = 12'b001010011010;
            14'b10_011000011110: DATA = 12'b001010011100;
            14'b10_011000011111: DATA = 12'b001010011110;
            14'b10_011000100000: DATA = 12'b001010100001;
            14'b10_011000100001: DATA = 12'b001010100011;
            14'b10_011000100010: DATA = 12'b001010100101;
            14'b10_011000100011: DATA = 12'b001010101000;
            14'b10_011000100100: DATA = 12'b001010101010;
            14'b10_011000100101: DATA = 12'b001010101100;
            14'b10_011000100110: DATA = 12'b001010101111;
            14'b10_011000100111: DATA = 12'b001010110001;
            14'b10_011000101000: DATA = 12'b001010110100;
            14'b10_011000101001: DATA = 12'b001010110110;
            14'b10_011000101010: DATA = 12'b001010111000;
            14'b10_011000101011: DATA = 12'b001010111011;
            14'b10_011000101100: DATA = 12'b001010111101;
            14'b10_011000101101: DATA = 12'b001010111111;
            14'b10_011000101110: DATA = 12'b001011000010;
            14'b10_011000101111: DATA = 12'b001011000100;
            14'b10_011000110000: DATA = 12'b001011000110;
            14'b10_011000110001: DATA = 12'b001011001001;
            14'b10_011000110010: DATA = 12'b001011001011;
            14'b10_011000110011: DATA = 12'b001011001110;
            14'b10_011000110100: DATA = 12'b001011010000;
            14'b10_011000110101: DATA = 12'b001011010010;
            14'b10_011000110110: DATA = 12'b001011010101;
            14'b10_011000110111: DATA = 12'b001011010111;
            14'b10_011000111000: DATA = 12'b001011011010;
            14'b10_011000111001: DATA = 12'b001011011100;
            14'b10_011000111010: DATA = 12'b001011011110;
            14'b10_011000111011: DATA = 12'b001011100001;
            14'b10_011000111100: DATA = 12'b001011100011;
            14'b10_011000111101: DATA = 12'b001011100110;
            14'b10_011000111110: DATA = 12'b001011101000;
            14'b10_011000111111: DATA = 12'b001011101010;
            14'b10_011001000000: DATA = 12'b001011101101;
            14'b10_011001000001: DATA = 12'b001011101111;
            14'b10_011001000010: DATA = 12'b001011110010;
            14'b10_011001000011: DATA = 12'b001011110100;
            14'b10_011001000100: DATA = 12'b001011110111;
            14'b10_011001000101: DATA = 12'b001011111001;
            14'b10_011001000110: DATA = 12'b001011111100;
            14'b10_011001000111: DATA = 12'b001011111110;
            14'b10_011001001000: DATA = 12'b001100000000;
            14'b10_011001001001: DATA = 12'b001100000011;
            14'b10_011001001010: DATA = 12'b001100000101;
            14'b10_011001001011: DATA = 12'b001100001000;
            14'b10_011001001100: DATA = 12'b001100001010;
            14'b10_011001001101: DATA = 12'b001100001101;
            14'b10_011001001110: DATA = 12'b001100001111;
            14'b10_011001001111: DATA = 12'b001100010010;
            14'b10_011001010000: DATA = 12'b001100010100;
            14'b10_011001010001: DATA = 12'b001100010111;
            14'b10_011001010010: DATA = 12'b001100011001;
            14'b10_011001010011: DATA = 12'b001100011100;
            14'b10_011001010100: DATA = 12'b001100011110;
            14'b10_011001010101: DATA = 12'b001100100001;
            14'b10_011001010110: DATA = 12'b001100100011;
            14'b10_011001010111: DATA = 12'b001100100110;
            14'b10_011001011000: DATA = 12'b001100101000;
            14'b10_011001011001: DATA = 12'b001100101011;
            14'b10_011001011010: DATA = 12'b001100101101;
            14'b10_011001011011: DATA = 12'b001100110000;
            14'b10_011001011100: DATA = 12'b001100110010;
            14'b10_011001011101: DATA = 12'b001100110101;
            14'b10_011001011110: DATA = 12'b001100110111;
            14'b10_011001011111: DATA = 12'b001100111010;
            14'b10_011001100000: DATA = 12'b001100111100;
            14'b10_011001100001: DATA = 12'b001100111111;
            14'b10_011001100010: DATA = 12'b001101000001;
            14'b10_011001100011: DATA = 12'b001101000100;
            14'b10_011001100100: DATA = 12'b001101000110;
            14'b10_011001100101: DATA = 12'b001101001001;
            14'b10_011001100110: DATA = 12'b001101001011;
            14'b10_011001100111: DATA = 12'b001101001110;
            14'b10_011001101000: DATA = 12'b001101010000;
            14'b10_011001101001: DATA = 12'b001101010011;
            14'b10_011001101010: DATA = 12'b001101010101;
            14'b10_011001101011: DATA = 12'b001101011000;
            14'b10_011001101100: DATA = 12'b001101011011;
            14'b10_011001101101: DATA = 12'b001101011101;
            14'b10_011001101110: DATA = 12'b001101100000;
            14'b10_011001101111: DATA = 12'b001101100010;
            14'b10_011001110000: DATA = 12'b001101100101;
            14'b10_011001110001: DATA = 12'b001101100111;
            14'b10_011001110010: DATA = 12'b001101101010;
            14'b10_011001110011: DATA = 12'b001101101101;
            14'b10_011001110100: DATA = 12'b001101101111;
            14'b10_011001110101: DATA = 12'b001101110010;
            14'b10_011001110110: DATA = 12'b001101110100;
            14'b10_011001110111: DATA = 12'b001101110111;
            14'b10_011001111000: DATA = 12'b001101111001;
            14'b10_011001111001: DATA = 12'b001101111100;
            14'b10_011001111010: DATA = 12'b001101111111;
            14'b10_011001111011: DATA = 12'b001110000001;
            14'b10_011001111100: DATA = 12'b001110000100;
            14'b10_011001111101: DATA = 12'b001110000110;
            14'b10_011001111110: DATA = 12'b001110001001;
            14'b10_011001111111: DATA = 12'b001110001100;
            14'b10_011010000000: DATA = 12'b001110001110;
            14'b10_011010000001: DATA = 12'b001110010001;
            14'b10_011010000010: DATA = 12'b001110010011;
            14'b10_011010000011: DATA = 12'b001110010110;
            14'b10_011010000100: DATA = 12'b001110011001;
            14'b10_011010000101: DATA = 12'b001110011011;
            14'b10_011010000110: DATA = 12'b001110011110;
            14'b10_011010000111: DATA = 12'b001110100001;
            14'b10_011010001000: DATA = 12'b001110100011;
            14'b10_011010001001: DATA = 12'b001110100110;
            14'b10_011010001010: DATA = 12'b001110101000;
            14'b10_011010001011: DATA = 12'b001110101011;
            14'b10_011010001100: DATA = 12'b001110101110;
            14'b10_011010001101: DATA = 12'b001110110000;
            14'b10_011010001110: DATA = 12'b001110110011;
            14'b10_011010001111: DATA = 12'b001110110110;
            14'b10_011010010000: DATA = 12'b001110111000;
            14'b10_011010010001: DATA = 12'b001110111011;
            14'b10_011010010010: DATA = 12'b001110111110;
            14'b10_011010010011: DATA = 12'b001111000000;
            14'b10_011010010100: DATA = 12'b001111000011;
            14'b10_011010010101: DATA = 12'b001111000110;
            14'b10_011010010110: DATA = 12'b001111001000;
            14'b10_011010010111: DATA = 12'b001111001011;
            14'b10_011010011000: DATA = 12'b001111001110;
            14'b10_011010011001: DATA = 12'b001111010000;
            14'b10_011010011010: DATA = 12'b001111010011;
            14'b10_011010011011: DATA = 12'b001111010110;
            14'b10_011010011100: DATA = 12'b001111011000;
            14'b10_011010011101: DATA = 12'b001111011011;
            14'b10_011010011110: DATA = 12'b001111011110;
            14'b10_011010011111: DATA = 12'b001111100000;
            14'b10_011010100000: DATA = 12'b001111100011;
            14'b10_011010100001: DATA = 12'b001111100110;
            14'b10_011010100010: DATA = 12'b001111101001;
            14'b10_011010100011: DATA = 12'b001111101011;
            14'b10_011010100100: DATA = 12'b001111101110;
            14'b10_011010100101: DATA = 12'b001111110001;
            14'b10_011010100110: DATA = 12'b001111110011;
            14'b10_011010100111: DATA = 12'b001111110110;
            14'b10_011010101000: DATA = 12'b001111111001;
            14'b10_011010101001: DATA = 12'b001111111011;
            14'b10_011010101010: DATA = 12'b001111111110;
            14'b10_011010101011: DATA = 12'b010000000001;
            14'b10_011010101100: DATA = 12'b010000000100;
            14'b10_011010101101: DATA = 12'b010000000110;
            14'b10_011010101110: DATA = 12'b010000001001;
            14'b10_011010101111: DATA = 12'b010000001100;
            14'b10_011010110000: DATA = 12'b010000001111;
            14'b10_011010110001: DATA = 12'b010000010001;
            14'b10_011010110010: DATA = 12'b010000010100;
            14'b10_011010110011: DATA = 12'b010000010111;
            14'b10_011010110100: DATA = 12'b010000011001;
            14'b10_011010110101: DATA = 12'b010000011100;
            14'b10_011010110110: DATA = 12'b010000011111;
            14'b10_011010110111: DATA = 12'b010000100010;
            14'b10_011010111000: DATA = 12'b010000100100;
            14'b10_011010111001: DATA = 12'b010000100111;
            14'b10_011010111010: DATA = 12'b010000101010;
            14'b10_011010111011: DATA = 12'b010000101101;
            14'b10_011010111100: DATA = 12'b010000101111;
            14'b10_011010111101: DATA = 12'b010000110010;
            14'b10_011010111110: DATA = 12'b010000110101;
            14'b10_011010111111: DATA = 12'b010000111000;
            14'b10_011011000000: DATA = 12'b010000111011;
            14'b10_011011000001: DATA = 12'b010000111101;
            14'b10_011011000010: DATA = 12'b010001000000;
            14'b10_011011000011: DATA = 12'b010001000011;
            14'b10_011011000100: DATA = 12'b010001000110;
            14'b10_011011000101: DATA = 12'b010001001000;
            14'b10_011011000110: DATA = 12'b010001001011;
            14'b10_011011000111: DATA = 12'b010001001110;
            14'b10_011011001000: DATA = 12'b010001010001;
            14'b10_011011001001: DATA = 12'b010001010100;
            14'b10_011011001010: DATA = 12'b010001010110;
            14'b10_011011001011: DATA = 12'b010001011001;
            14'b10_011011001100: DATA = 12'b010001011100;
            14'b10_011011001101: DATA = 12'b010001011111;
            14'b10_011011001110: DATA = 12'b010001100010;
            14'b10_011011001111: DATA = 12'b010001100100;
            14'b10_011011010000: DATA = 12'b010001100111;
            14'b10_011011010001: DATA = 12'b010001101010;
            14'b10_011011010010: DATA = 12'b010001101101;
            14'b10_011011010011: DATA = 12'b010001110000;
            14'b10_011011010100: DATA = 12'b010001110010;
            14'b10_011011010101: DATA = 12'b010001110101;
            14'b10_011011010110: DATA = 12'b010001111000;
            14'b10_011011010111: DATA = 12'b010001111011;
            14'b10_011011011000: DATA = 12'b010001111110;
            14'b10_011011011001: DATA = 12'b010010000000;
            14'b10_011011011010: DATA = 12'b010010000011;
            14'b10_011011011011: DATA = 12'b010010000110;
            14'b10_011011011100: DATA = 12'b010010001001;
            14'b10_011011011101: DATA = 12'b010010001100;
            14'b10_011011011110: DATA = 12'b010010001111;
            14'b10_011011011111: DATA = 12'b010010010001;
            14'b10_011011100000: DATA = 12'b010010010100;
            14'b10_011011100001: DATA = 12'b010010010111;
            14'b10_011011100010: DATA = 12'b010010011010;
            14'b10_011011100011: DATA = 12'b010010011101;
            14'b10_011011100100: DATA = 12'b010010100000;
            14'b10_011011100101: DATA = 12'b010010100011;
            14'b10_011011100110: DATA = 12'b010010100101;
            14'b10_011011100111: DATA = 12'b010010101000;
            14'b10_011011101000: DATA = 12'b010010101011;
            14'b10_011011101001: DATA = 12'b010010101110;
            14'b10_011011101010: DATA = 12'b010010110001;
            14'b10_011011101011: DATA = 12'b010010110100;
            14'b10_011011101100: DATA = 12'b010010110111;
            14'b10_011011101101: DATA = 12'b010010111001;
            14'b10_011011101110: DATA = 12'b010010111100;
            14'b10_011011101111: DATA = 12'b010010111111;
            14'b10_011011110000: DATA = 12'b010011000010;
            14'b10_011011110001: DATA = 12'b010011000101;
            14'b10_011011110010: DATA = 12'b010011001000;
            14'b10_011011110011: DATA = 12'b010011001011;
            14'b10_011011110100: DATA = 12'b010011001101;
            14'b10_011011110101: DATA = 12'b010011010000;
            14'b10_011011110110: DATA = 12'b010011010011;
            14'b10_011011110111: DATA = 12'b010011010110;
            14'b10_011011111000: DATA = 12'b010011011001;
            14'b10_011011111001: DATA = 12'b010011011100;
            14'b10_011011111010: DATA = 12'b010011011111;
            14'b10_011011111011: DATA = 12'b010011100010;
            14'b10_011011111100: DATA = 12'b010011100101;
            14'b10_011011111101: DATA = 12'b010011100111;
            14'b10_011011111110: DATA = 12'b010011101010;
            14'b10_011011111111: DATA = 12'b010011101101;
            14'b10_011100000000: DATA = 12'b010011110000;
            14'b10_011100000001: DATA = 12'b010011110011;
            14'b10_011100000010: DATA = 12'b010011110110;
            14'b10_011100000011: DATA = 12'b010011111001;
            14'b10_011100000100: DATA = 12'b010011111100;
            14'b10_011100000101: DATA = 12'b010011111111;
            14'b10_011100000110: DATA = 12'b010100000010;
            14'b10_011100000111: DATA = 12'b010100000100;
            14'b10_011100001000: DATA = 12'b010100000111;
            14'b10_011100001001: DATA = 12'b010100001010;
            14'b10_011100001010: DATA = 12'b010100001101;
            14'b10_011100001011: DATA = 12'b010100010000;
            14'b10_011100001100: DATA = 12'b010100010011;
            14'b10_011100001101: DATA = 12'b010100010110;
            14'b10_011100001110: DATA = 12'b010100011001;
            14'b10_011100001111: DATA = 12'b010100011100;
            14'b10_011100010000: DATA = 12'b010100011111;
            14'b10_011100010001: DATA = 12'b010100100010;
            14'b10_011100010010: DATA = 12'b010100100101;
            14'b10_011100010011: DATA = 12'b010100101000;
            14'b10_011100010100: DATA = 12'b010100101011;
            14'b10_011100010101: DATA = 12'b010100101101;
            14'b10_011100010110: DATA = 12'b010100110000;
            14'b10_011100010111: DATA = 12'b010100110011;
            14'b10_011100011000: DATA = 12'b010100110110;
            14'b10_011100011001: DATA = 12'b010100111001;
            14'b10_011100011010: DATA = 12'b010100111100;
            14'b10_011100011011: DATA = 12'b010100111111;
            14'b10_011100011100: DATA = 12'b010101000010;
            14'b10_011100011101: DATA = 12'b010101000101;
            14'b10_011100011110: DATA = 12'b010101001000;
            14'b10_011100011111: DATA = 12'b010101001011;
            14'b10_011100100000: DATA = 12'b010101001110;
            14'b10_011100100001: DATA = 12'b010101010001;
            14'b10_011100100010: DATA = 12'b010101010100;
            14'b10_011100100011: DATA = 12'b010101010111;
            14'b10_011100100100: DATA = 12'b010101011010;
            14'b10_011100100101: DATA = 12'b010101011101;
            14'b10_011100100110: DATA = 12'b010101100000;
            14'b10_011100100111: DATA = 12'b010101100011;
            14'b10_011100101000: DATA = 12'b010101100110;
            14'b10_011100101001: DATA = 12'b010101101001;
            14'b10_011100101010: DATA = 12'b010101101100;
            14'b10_011100101011: DATA = 12'b010101101111;
            14'b10_011100101100: DATA = 12'b010101110001;
            14'b10_011100101101: DATA = 12'b010101110100;
            14'b10_011100101110: DATA = 12'b010101110111;
            14'b10_011100101111: DATA = 12'b010101111010;
            14'b10_011100110000: DATA = 12'b010101111101;
            14'b10_011100110001: DATA = 12'b010110000000;
            14'b10_011100110010: DATA = 12'b010110000011;
            14'b10_011100110011: DATA = 12'b010110000110;
            14'b10_011100110100: DATA = 12'b010110001001;
            14'b10_011100110101: DATA = 12'b010110001100;
            14'b10_011100110110: DATA = 12'b010110001111;
            14'b10_011100110111: DATA = 12'b010110010010;
            14'b10_011100111000: DATA = 12'b010110010101;
            14'b10_011100111001: DATA = 12'b010110011000;
            14'b10_011100111010: DATA = 12'b010110011011;
            14'b10_011100111011: DATA = 12'b010110011110;
            14'b10_011100111100: DATA = 12'b010110100001;
            14'b10_011100111101: DATA = 12'b010110100100;
            14'b10_011100111110: DATA = 12'b010110100111;
            14'b10_011100111111: DATA = 12'b010110101010;
            14'b10_011101000000: DATA = 12'b010110101101;
            14'b10_011101000001: DATA = 12'b010110110000;
            14'b10_011101000010: DATA = 12'b010110110011;
            14'b10_011101000011: DATA = 12'b010110110110;
            14'b10_011101000100: DATA = 12'b010110111001;
            14'b10_011101000101: DATA = 12'b010110111100;
            14'b10_011101000110: DATA = 12'b010110111111;
            14'b10_011101000111: DATA = 12'b010111000010;
            14'b10_011101001000: DATA = 12'b010111000101;
            14'b10_011101001001: DATA = 12'b010111001000;
            14'b10_011101001010: DATA = 12'b010111001011;
            14'b10_011101001011: DATA = 12'b010111001110;
            14'b10_011101001100: DATA = 12'b010111010001;
            14'b10_011101001101: DATA = 12'b010111010100;
            14'b10_011101001110: DATA = 12'b010111010111;
            14'b10_011101001111: DATA = 12'b010111011011;
            14'b10_011101010000: DATA = 12'b010111011110;
            14'b10_011101010001: DATA = 12'b010111100001;
            14'b10_011101010010: DATA = 12'b010111100100;
            14'b10_011101010011: DATA = 12'b010111100111;
            14'b10_011101010100: DATA = 12'b010111101010;
            14'b10_011101010101: DATA = 12'b010111101101;
            14'b10_011101010110: DATA = 12'b010111110000;
            14'b10_011101010111: DATA = 12'b010111110011;
            14'b10_011101011000: DATA = 12'b010111110110;
            14'b10_011101011001: DATA = 12'b010111111001;
            14'b10_011101011010: DATA = 12'b010111111100;
            14'b10_011101011011: DATA = 12'b010111111111;
            14'b10_011101011100: DATA = 12'b011000000010;
            14'b10_011101011101: DATA = 12'b011000000101;
            14'b10_011101011110: DATA = 12'b011000001000;
            14'b10_011101011111: DATA = 12'b011000001011;
            14'b10_011101100000: DATA = 12'b011000001110;
            14'b10_011101100001: DATA = 12'b011000010001;
            14'b10_011101100010: DATA = 12'b011000010100;
            14'b10_011101100011: DATA = 12'b011000010111;
            14'b10_011101100100: DATA = 12'b011000011010;
            14'b10_011101100101: DATA = 12'b011000011101;
            14'b10_011101100110: DATA = 12'b011000100000;
            14'b10_011101100111: DATA = 12'b011000100011;
            14'b10_011101101000: DATA = 12'b011000100111;
            14'b10_011101101001: DATA = 12'b011000101010;
            14'b10_011101101010: DATA = 12'b011000101101;
            14'b10_011101101011: DATA = 12'b011000110000;
            14'b10_011101101100: DATA = 12'b011000110011;
            14'b10_011101101101: DATA = 12'b011000110110;
            14'b10_011101101110: DATA = 12'b011000111001;
            14'b10_011101101111: DATA = 12'b011000111100;
            14'b10_011101110000: DATA = 12'b011000111111;
            14'b10_011101110001: DATA = 12'b011001000010;
            14'b10_011101110010: DATA = 12'b011001000101;
            14'b10_011101110011: DATA = 12'b011001001000;
            14'b10_011101110100: DATA = 12'b011001001011;
            14'b10_011101110101: DATA = 12'b011001001110;
            14'b10_011101110110: DATA = 12'b011001010001;
            14'b10_011101110111: DATA = 12'b011001010100;
            14'b10_011101111000: DATA = 12'b011001011000;
            14'b10_011101111001: DATA = 12'b011001011011;
            14'b10_011101111010: DATA = 12'b011001011110;
            14'b10_011101111011: DATA = 12'b011001100001;
            14'b10_011101111100: DATA = 12'b011001100100;
            14'b10_011101111101: DATA = 12'b011001100111;
            14'b10_011101111110: DATA = 12'b011001101010;
            14'b10_011101111111: DATA = 12'b011001101101;
            14'b10_011110000000: DATA = 12'b011001110000;
            14'b10_011110000001: DATA = 12'b011001110011;
            14'b10_011110000010: DATA = 12'b011001110110;
            14'b10_011110000011: DATA = 12'b011001111001;
            14'b10_011110000100: DATA = 12'b011001111100;
            14'b10_011110000101: DATA = 12'b011010000000;
            14'b10_011110000110: DATA = 12'b011010000011;
            14'b10_011110000111: DATA = 12'b011010000110;
            14'b10_011110001000: DATA = 12'b011010001001;
            14'b10_011110001001: DATA = 12'b011010001100;
            14'b10_011110001010: DATA = 12'b011010001111;
            14'b10_011110001011: DATA = 12'b011010010010;
            14'b10_011110001100: DATA = 12'b011010010101;
            14'b10_011110001101: DATA = 12'b011010011000;
            14'b10_011110001110: DATA = 12'b011010011011;
            14'b10_011110001111: DATA = 12'b011010011110;
            14'b10_011110010000: DATA = 12'b011010100010;
            14'b10_011110010001: DATA = 12'b011010100101;
            14'b10_011110010010: DATA = 12'b011010101000;
            14'b10_011110010011: DATA = 12'b011010101011;
            14'b10_011110010100: DATA = 12'b011010101110;
            14'b10_011110010101: DATA = 12'b011010110001;
            14'b10_011110010110: DATA = 12'b011010110100;
            14'b10_011110010111: DATA = 12'b011010110111;
            14'b10_011110011000: DATA = 12'b011010111010;
            14'b10_011110011001: DATA = 12'b011010111101;
            14'b10_011110011010: DATA = 12'b011011000001;
            14'b10_011110011011: DATA = 12'b011011000100;
            14'b10_011110011100: DATA = 12'b011011000111;
            14'b10_011110011101: DATA = 12'b011011001010;
            14'b10_011110011110: DATA = 12'b011011001101;
            14'b10_011110011111: DATA = 12'b011011010000;
            14'b10_011110100000: DATA = 12'b011011010011;
            14'b10_011110100001: DATA = 12'b011011010110;
            14'b10_011110100010: DATA = 12'b011011011001;
            14'b10_011110100011: DATA = 12'b011011011100;
            14'b10_011110100100: DATA = 12'b011011100000;
            14'b10_011110100101: DATA = 12'b011011100011;
            14'b10_011110100110: DATA = 12'b011011100110;
            14'b10_011110100111: DATA = 12'b011011101001;
            14'b10_011110101000: DATA = 12'b011011101100;
            14'b10_011110101001: DATA = 12'b011011101111;
            14'b10_011110101010: DATA = 12'b011011110010;
            14'b10_011110101011: DATA = 12'b011011110101;
            14'b10_011110101100: DATA = 12'b011011111000;
            14'b10_011110101101: DATA = 12'b011011111100;
            14'b10_011110101110: DATA = 12'b011011111111;
            14'b10_011110101111: DATA = 12'b011100000010;
            14'b10_011110110000: DATA = 12'b011100000101;
            14'b10_011110110001: DATA = 12'b011100001000;
            14'b10_011110110010: DATA = 12'b011100001011;
            14'b10_011110110011: DATA = 12'b011100001110;
            14'b10_011110110100: DATA = 12'b011100010001;
            14'b10_011110110101: DATA = 12'b011100010101;
            14'b10_011110110110: DATA = 12'b011100011000;
            14'b10_011110110111: DATA = 12'b011100011011;
            14'b10_011110111000: DATA = 12'b011100011110;
            14'b10_011110111001: DATA = 12'b011100100001;
            14'b10_011110111010: DATA = 12'b011100100100;
            14'b10_011110111011: DATA = 12'b011100100111;
            14'b10_011110111100: DATA = 12'b011100101010;
            14'b10_011110111101: DATA = 12'b011100101101;
            14'b10_011110111110: DATA = 12'b011100110001;
            14'b10_011110111111: DATA = 12'b011100110100;
            14'b10_011111000000: DATA = 12'b011100110111;
            14'b10_011111000001: DATA = 12'b011100111010;
            14'b10_011111000010: DATA = 12'b011100111101;
            14'b10_011111000011: DATA = 12'b011101000000;
            14'b10_011111000100: DATA = 12'b011101000011;
            14'b10_011111000101: DATA = 12'b011101000110;
            14'b10_011111000110: DATA = 12'b011101001010;
            14'b10_011111000111: DATA = 12'b011101001101;
            14'b10_011111001000: DATA = 12'b011101010000;
            14'b10_011111001001: DATA = 12'b011101010011;
            14'b10_011111001010: DATA = 12'b011101010110;
            14'b10_011111001011: DATA = 12'b011101011001;
            14'b10_011111001100: DATA = 12'b011101011100;
            14'b10_011111001101: DATA = 12'b011101100000;
            14'b10_011111001110: DATA = 12'b011101100011;
            14'b10_011111001111: DATA = 12'b011101100110;
            14'b10_011111010000: DATA = 12'b011101101001;
            14'b10_011111010001: DATA = 12'b011101101100;
            14'b10_011111010010: DATA = 12'b011101101111;
            14'b10_011111010011: DATA = 12'b011101110010;
            14'b10_011111010100: DATA = 12'b011101110101;
            14'b10_011111010101: DATA = 12'b011101111001;
            14'b10_011111010110: DATA = 12'b011101111100;
            14'b10_011111010111: DATA = 12'b011101111111;
            14'b10_011111011000: DATA = 12'b011110000010;
            14'b10_011111011001: DATA = 12'b011110000101;
            14'b10_011111011010: DATA = 12'b011110001000;
            14'b10_011111011011: DATA = 12'b011110001011;
            14'b10_011111011100: DATA = 12'b011110001111;
            14'b10_011111011101: DATA = 12'b011110010010;
            14'b10_011111011110: DATA = 12'b011110010101;
            14'b10_011111011111: DATA = 12'b011110011000;
            14'b10_011111100000: DATA = 12'b011110011011;
            14'b10_011111100001: DATA = 12'b011110011110;
            14'b10_011111100010: DATA = 12'b011110100001;
            14'b10_011111100011: DATA = 12'b011110100100;
            14'b10_011111100100: DATA = 12'b011110101000;
            14'b10_011111100101: DATA = 12'b011110101011;
            14'b10_011111100110: DATA = 12'b011110101110;
            14'b10_011111100111: DATA = 12'b011110110001;
            14'b10_011111101000: DATA = 12'b011110110100;
            14'b10_011111101001: DATA = 12'b011110110111;
            14'b10_011111101010: DATA = 12'b011110111010;
            14'b10_011111101011: DATA = 12'b011110111110;
            14'b10_011111101100: DATA = 12'b011111000001;
            14'b10_011111101101: DATA = 12'b011111000100;
            14'b10_011111101110: DATA = 12'b011111000111;
            14'b10_011111101111: DATA = 12'b011111001010;
            14'b10_011111110000: DATA = 12'b011111001101;
            14'b10_011111110001: DATA = 12'b011111010000;
            14'b10_011111110010: DATA = 12'b011111010100;
            14'b10_011111110011: DATA = 12'b011111010111;
            14'b10_011111110100: DATA = 12'b011111011010;
            14'b10_011111110101: DATA = 12'b011111011101;
            14'b10_011111110110: DATA = 12'b011111100000;
            14'b10_011111110111: DATA = 12'b011111100011;
            14'b10_011111111000: DATA = 12'b011111100110;
            14'b10_011111111001: DATA = 12'b011111101010;
            14'b10_011111111010: DATA = 12'b011111101101;
            14'b10_011111111011: DATA = 12'b011111110000;
            14'b10_011111111100: DATA = 12'b011111110011;
            14'b10_011111111101: DATA = 12'b011111110110;
            14'b10_011111111110: DATA = 12'b011111111001;
            14'b10_011111111111: DATA = 12'b011111111100;
            14'b10_100000000000: DATA = 12'b011111111111;
            14'b10_100000000001: DATA = 12'b100000000011;
            14'b10_100000000010: DATA = 12'b100000000110;
            14'b10_100000000011: DATA = 12'b100000001001;
            14'b10_100000000100: DATA = 12'b100000001100;
            14'b10_100000000101: DATA = 12'b100000001111;
            14'b10_100000000110: DATA = 12'b100000010010;
            14'b10_100000000111: DATA = 12'b100000010101;
            14'b10_100000001000: DATA = 12'b100000011001;
            14'b10_100000001001: DATA = 12'b100000011100;
            14'b10_100000001010: DATA = 12'b100000011111;
            14'b10_100000001011: DATA = 12'b100000100010;
            14'b10_100000001100: DATA = 12'b100000100101;
            14'b10_100000001101: DATA = 12'b100000101000;
            14'b10_100000001110: DATA = 12'b100000101011;
            14'b10_100000001111: DATA = 12'b100000101111;
            14'b10_100000010000: DATA = 12'b100000110010;
            14'b10_100000010001: DATA = 12'b100000110101;
            14'b10_100000010010: DATA = 12'b100000111000;
            14'b10_100000010011: DATA = 12'b100000111011;
            14'b10_100000010100: DATA = 12'b100000111110;
            14'b10_100000010101: DATA = 12'b100001000001;
            14'b10_100000010110: DATA = 12'b100001000101;
            14'b10_100000010111: DATA = 12'b100001001000;
            14'b10_100000011000: DATA = 12'b100001001011;
            14'b10_100000011001: DATA = 12'b100001001110;
            14'b10_100000011010: DATA = 12'b100001010001;
            14'b10_100000011011: DATA = 12'b100001010100;
            14'b10_100000011100: DATA = 12'b100001010111;
            14'b10_100000011101: DATA = 12'b100001011011;
            14'b10_100000011110: DATA = 12'b100001011110;
            14'b10_100000011111: DATA = 12'b100001100001;
            14'b10_100000100000: DATA = 12'b100001100100;
            14'b10_100000100001: DATA = 12'b100001100111;
            14'b10_100000100010: DATA = 12'b100001101010;
            14'b10_100000100011: DATA = 12'b100001101101;
            14'b10_100000100100: DATA = 12'b100001110000;
            14'b10_100000100101: DATA = 12'b100001110100;
            14'b10_100000100110: DATA = 12'b100001110111;
            14'b10_100000100111: DATA = 12'b100001111010;
            14'b10_100000101000: DATA = 12'b100001111101;
            14'b10_100000101001: DATA = 12'b100010000000;
            14'b10_100000101010: DATA = 12'b100010000011;
            14'b10_100000101011: DATA = 12'b100010000110;
            14'b10_100000101100: DATA = 12'b100010001010;
            14'b10_100000101101: DATA = 12'b100010001101;
            14'b10_100000101110: DATA = 12'b100010010000;
            14'b10_100000101111: DATA = 12'b100010010011;
            14'b10_100000110000: DATA = 12'b100010010110;
            14'b10_100000110001: DATA = 12'b100010011001;
            14'b10_100000110010: DATA = 12'b100010011100;
            14'b10_100000110011: DATA = 12'b100010011111;
            14'b10_100000110100: DATA = 12'b100010100011;
            14'b10_100000110101: DATA = 12'b100010100110;
            14'b10_100000110110: DATA = 12'b100010101001;
            14'b10_100000110111: DATA = 12'b100010101100;
            14'b10_100000111000: DATA = 12'b100010101111;
            14'b10_100000111001: DATA = 12'b100010110010;
            14'b10_100000111010: DATA = 12'b100010110101;
            14'b10_100000111011: DATA = 12'b100010111001;
            14'b10_100000111100: DATA = 12'b100010111100;
            14'b10_100000111101: DATA = 12'b100010111111;
            14'b10_100000111110: DATA = 12'b100011000010;
            14'b10_100000111111: DATA = 12'b100011000101;
            14'b10_100001000000: DATA = 12'b100011001000;
            14'b10_100001000001: DATA = 12'b100011001011;
            14'b10_100001000010: DATA = 12'b100011001110;
            14'b10_100001000011: DATA = 12'b100011010010;
            14'b10_100001000100: DATA = 12'b100011010101;
            14'b10_100001000101: DATA = 12'b100011011000;
            14'b10_100001000110: DATA = 12'b100011011011;
            14'b10_100001000111: DATA = 12'b100011011110;
            14'b10_100001001000: DATA = 12'b100011100001;
            14'b10_100001001001: DATA = 12'b100011100100;
            14'b10_100001001010: DATA = 12'b100011100111;
            14'b10_100001001011: DATA = 12'b100011101010;
            14'b10_100001001100: DATA = 12'b100011101110;
            14'b10_100001001101: DATA = 12'b100011110001;
            14'b10_100001001110: DATA = 12'b100011110100;
            14'b10_100001001111: DATA = 12'b100011110111;
            14'b10_100001010000: DATA = 12'b100011111010;
            14'b10_100001010001: DATA = 12'b100011111101;
            14'b10_100001010010: DATA = 12'b100100000000;
            14'b10_100001010011: DATA = 12'b100100000011;
            14'b10_100001010100: DATA = 12'b100100000111;
            14'b10_100001010101: DATA = 12'b100100001010;
            14'b10_100001010110: DATA = 12'b100100001101;
            14'b10_100001010111: DATA = 12'b100100010000;
            14'b10_100001011000: DATA = 12'b100100010011;
            14'b10_100001011001: DATA = 12'b100100010110;
            14'b10_100001011010: DATA = 12'b100100011001;
            14'b10_100001011011: DATA = 12'b100100011100;
            14'b10_100001011100: DATA = 12'b100100011111;
            14'b10_100001011101: DATA = 12'b100100100011;
            14'b10_100001011110: DATA = 12'b100100100110;
            14'b10_100001011111: DATA = 12'b100100101001;
            14'b10_100001100000: DATA = 12'b100100101100;
            14'b10_100001100001: DATA = 12'b100100101111;
            14'b10_100001100010: DATA = 12'b100100110010;
            14'b10_100001100011: DATA = 12'b100100110101;
            14'b10_100001100100: DATA = 12'b100100111000;
            14'b10_100001100101: DATA = 12'b100100111011;
            14'b10_100001100110: DATA = 12'b100100111110;
            14'b10_100001100111: DATA = 12'b100101000010;
            14'b10_100001101000: DATA = 12'b100101000101;
            14'b10_100001101001: DATA = 12'b100101001000;
            14'b10_100001101010: DATA = 12'b100101001011;
            14'b10_100001101011: DATA = 12'b100101001110;
            14'b10_100001101100: DATA = 12'b100101010001;
            14'b10_100001101101: DATA = 12'b100101010100;
            14'b10_100001101110: DATA = 12'b100101010111;
            14'b10_100001101111: DATA = 12'b100101011010;
            14'b10_100001110000: DATA = 12'b100101011101;
            14'b10_100001110001: DATA = 12'b100101100001;
            14'b10_100001110010: DATA = 12'b100101100100;
            14'b10_100001110011: DATA = 12'b100101100111;
            14'b10_100001110100: DATA = 12'b100101101010;
            14'b10_100001110101: DATA = 12'b100101101101;
            14'b10_100001110110: DATA = 12'b100101110000;
            14'b10_100001110111: DATA = 12'b100101110011;
            14'b10_100001111000: DATA = 12'b100101110110;
            14'b10_100001111001: DATA = 12'b100101111001;
            14'b10_100001111010: DATA = 12'b100101111100;
            14'b10_100001111011: DATA = 12'b100101111111;
            14'b10_100001111100: DATA = 12'b100110000011;
            14'b10_100001111101: DATA = 12'b100110000110;
            14'b10_100001111110: DATA = 12'b100110001001;
            14'b10_100001111111: DATA = 12'b100110001100;
            14'b10_100010000000: DATA = 12'b100110001111;
            14'b10_100010000001: DATA = 12'b100110010010;
            14'b10_100010000010: DATA = 12'b100110010101;
            14'b10_100010000011: DATA = 12'b100110011000;
            14'b10_100010000100: DATA = 12'b100110011011;
            14'b10_100010000101: DATA = 12'b100110011110;
            14'b10_100010000110: DATA = 12'b100110100001;
            14'b10_100010000111: DATA = 12'b100110100100;
            14'b10_100010001000: DATA = 12'b100110100111;
            14'b10_100010001001: DATA = 12'b100110101011;
            14'b10_100010001010: DATA = 12'b100110101110;
            14'b10_100010001011: DATA = 12'b100110110001;
            14'b10_100010001100: DATA = 12'b100110110100;
            14'b10_100010001101: DATA = 12'b100110110111;
            14'b10_100010001110: DATA = 12'b100110111010;
            14'b10_100010001111: DATA = 12'b100110111101;
            14'b10_100010010000: DATA = 12'b100111000000;
            14'b10_100010010001: DATA = 12'b100111000011;
            14'b10_100010010010: DATA = 12'b100111000110;
            14'b10_100010010011: DATA = 12'b100111001001;
            14'b10_100010010100: DATA = 12'b100111001100;
            14'b10_100010010101: DATA = 12'b100111001111;
            14'b10_100010010110: DATA = 12'b100111010010;
            14'b10_100010010111: DATA = 12'b100111010101;
            14'b10_100010011000: DATA = 12'b100111011000;
            14'b10_100010011001: DATA = 12'b100111011100;
            14'b10_100010011010: DATA = 12'b100111011111;
            14'b10_100010011011: DATA = 12'b100111100010;
            14'b10_100010011100: DATA = 12'b100111100101;
            14'b10_100010011101: DATA = 12'b100111101000;
            14'b10_100010011110: DATA = 12'b100111101011;
            14'b10_100010011111: DATA = 12'b100111101110;
            14'b10_100010100000: DATA = 12'b100111110001;
            14'b10_100010100001: DATA = 12'b100111110100;
            14'b10_100010100010: DATA = 12'b100111110111;
            14'b10_100010100011: DATA = 12'b100111111010;
            14'b10_100010100100: DATA = 12'b100111111101;
            14'b10_100010100101: DATA = 12'b101000000000;
            14'b10_100010100110: DATA = 12'b101000000011;
            14'b10_100010100111: DATA = 12'b101000000110;
            14'b10_100010101000: DATA = 12'b101000001001;
            14'b10_100010101001: DATA = 12'b101000001100;
            14'b10_100010101010: DATA = 12'b101000001111;
            14'b10_100010101011: DATA = 12'b101000010010;
            14'b10_100010101100: DATA = 12'b101000010101;
            14'b10_100010101101: DATA = 12'b101000011000;
            14'b10_100010101110: DATA = 12'b101000011011;
            14'b10_100010101111: DATA = 12'b101000011110;
            14'b10_100010110000: DATA = 12'b101000100001;
            14'b10_100010110001: DATA = 12'b101000100100;
            14'b10_100010110010: DATA = 12'b101000101000;
            14'b10_100010110011: DATA = 12'b101000101011;
            14'b10_100010110100: DATA = 12'b101000101110;
            14'b10_100010110101: DATA = 12'b101000110001;
            14'b10_100010110110: DATA = 12'b101000110100;
            14'b10_100010110111: DATA = 12'b101000110111;
            14'b10_100010111000: DATA = 12'b101000111010;
            14'b10_100010111001: DATA = 12'b101000111101;
            14'b10_100010111010: DATA = 12'b101001000000;
            14'b10_100010111011: DATA = 12'b101001000011;
            14'b10_100010111100: DATA = 12'b101001000110;
            14'b10_100010111101: DATA = 12'b101001001001;
            14'b10_100010111110: DATA = 12'b101001001100;
            14'b10_100010111111: DATA = 12'b101001001111;
            14'b10_100011000000: DATA = 12'b101001010010;
            14'b10_100011000001: DATA = 12'b101001010101;
            14'b10_100011000010: DATA = 12'b101001011000;
            14'b10_100011000011: DATA = 12'b101001011011;
            14'b10_100011000100: DATA = 12'b101001011110;
            14'b10_100011000101: DATA = 12'b101001100001;
            14'b10_100011000110: DATA = 12'b101001100100;
            14'b10_100011000111: DATA = 12'b101001100111;
            14'b10_100011001000: DATA = 12'b101001101010;
            14'b10_100011001001: DATA = 12'b101001101101;
            14'b10_100011001010: DATA = 12'b101001110000;
            14'b10_100011001011: DATA = 12'b101001110011;
            14'b10_100011001100: DATA = 12'b101001110110;
            14'b10_100011001101: DATA = 12'b101001111001;
            14'b10_100011001110: DATA = 12'b101001111100;
            14'b10_100011001111: DATA = 12'b101001111111;
            14'b10_100011010000: DATA = 12'b101010000010;
            14'b10_100011010001: DATA = 12'b101010000101;
            14'b10_100011010010: DATA = 12'b101010001000;
            14'b10_100011010011: DATA = 12'b101010001011;
            14'b10_100011010100: DATA = 12'b101010001110;
            14'b10_100011010101: DATA = 12'b101010010000;
            14'b10_100011010110: DATA = 12'b101010010011;
            14'b10_100011010111: DATA = 12'b101010010110;
            14'b10_100011011000: DATA = 12'b101010011001;
            14'b10_100011011001: DATA = 12'b101010011100;
            14'b10_100011011010: DATA = 12'b101010011111;
            14'b10_100011011011: DATA = 12'b101010100010;
            14'b10_100011011100: DATA = 12'b101010100101;
            14'b10_100011011101: DATA = 12'b101010101000;
            14'b10_100011011110: DATA = 12'b101010101011;
            14'b10_100011011111: DATA = 12'b101010101110;
            14'b10_100011100000: DATA = 12'b101010110001;
            14'b10_100011100001: DATA = 12'b101010110100;
            14'b10_100011100010: DATA = 12'b101010110111;
            14'b10_100011100011: DATA = 12'b101010111010;
            14'b10_100011100100: DATA = 12'b101010111101;
            14'b10_100011100101: DATA = 12'b101011000000;
            14'b10_100011100110: DATA = 12'b101011000011;
            14'b10_100011100111: DATA = 12'b101011000110;
            14'b10_100011101000: DATA = 12'b101011001001;
            14'b10_100011101001: DATA = 12'b101011001100;
            14'b10_100011101010: DATA = 12'b101011001111;
            14'b10_100011101011: DATA = 12'b101011010010;
            14'b10_100011101100: DATA = 12'b101011010100;
            14'b10_100011101101: DATA = 12'b101011010111;
            14'b10_100011101110: DATA = 12'b101011011010;
            14'b10_100011101111: DATA = 12'b101011011101;
            14'b10_100011110000: DATA = 12'b101011100000;
            14'b10_100011110001: DATA = 12'b101011100011;
            14'b10_100011110010: DATA = 12'b101011100110;
            14'b10_100011110011: DATA = 12'b101011101001;
            14'b10_100011110100: DATA = 12'b101011101100;
            14'b10_100011110101: DATA = 12'b101011101111;
            14'b10_100011110110: DATA = 12'b101011110010;
            14'b10_100011110111: DATA = 12'b101011110101;
            14'b10_100011111000: DATA = 12'b101011111000;
            14'b10_100011111001: DATA = 12'b101011111011;
            14'b10_100011111010: DATA = 12'b101011111101;
            14'b10_100011111011: DATA = 12'b101100000000;
            14'b10_100011111100: DATA = 12'b101100000011;
            14'b10_100011111101: DATA = 12'b101100000110;
            14'b10_100011111110: DATA = 12'b101100001001;
            14'b10_100011111111: DATA = 12'b101100001100;
            14'b10_100100000000: DATA = 12'b101100001111;
            14'b10_100100000001: DATA = 12'b101100010010;
            14'b10_100100000010: DATA = 12'b101100010101;
            14'b10_100100000011: DATA = 12'b101100011000;
            14'b10_100100000100: DATA = 12'b101100011010;
            14'b10_100100000101: DATA = 12'b101100011101;
            14'b10_100100000110: DATA = 12'b101100100000;
            14'b10_100100000111: DATA = 12'b101100100011;
            14'b10_100100001000: DATA = 12'b101100100110;
            14'b10_100100001001: DATA = 12'b101100101001;
            14'b10_100100001010: DATA = 12'b101100101100;
            14'b10_100100001011: DATA = 12'b101100101111;
            14'b10_100100001100: DATA = 12'b101100110010;
            14'b10_100100001101: DATA = 12'b101100110100;
            14'b10_100100001110: DATA = 12'b101100110111;
            14'b10_100100001111: DATA = 12'b101100111010;
            14'b10_100100010000: DATA = 12'b101100111101;
            14'b10_100100010001: DATA = 12'b101101000000;
            14'b10_100100010010: DATA = 12'b101101000011;
            14'b10_100100010011: DATA = 12'b101101000110;
            14'b10_100100010100: DATA = 12'b101101001000;
            14'b10_100100010101: DATA = 12'b101101001011;
            14'b10_100100010110: DATA = 12'b101101001110;
            14'b10_100100010111: DATA = 12'b101101010001;
            14'b10_100100011000: DATA = 12'b101101010100;
            14'b10_100100011001: DATA = 12'b101101010111;
            14'b10_100100011010: DATA = 12'b101101011010;
            14'b10_100100011011: DATA = 12'b101101011100;
            14'b10_100100011100: DATA = 12'b101101011111;
            14'b10_100100011101: DATA = 12'b101101100010;
            14'b10_100100011110: DATA = 12'b101101100101;
            14'b10_100100011111: DATA = 12'b101101101000;
            14'b10_100100100000: DATA = 12'b101101101011;
            14'b10_100100100001: DATA = 12'b101101101110;
            14'b10_100100100010: DATA = 12'b101101110000;
            14'b10_100100100011: DATA = 12'b101101110011;
            14'b10_100100100100: DATA = 12'b101101110110;
            14'b10_100100100101: DATA = 12'b101101111001;
            14'b10_100100100110: DATA = 12'b101101111100;
            14'b10_100100100111: DATA = 12'b101101111111;
            14'b10_100100101000: DATA = 12'b101110000001;
            14'b10_100100101001: DATA = 12'b101110000100;
            14'b10_100100101010: DATA = 12'b101110000111;
            14'b10_100100101011: DATA = 12'b101110001010;
            14'b10_100100101100: DATA = 12'b101110001101;
            14'b10_100100101101: DATA = 12'b101110001111;
            14'b10_100100101110: DATA = 12'b101110010010;
            14'b10_100100101111: DATA = 12'b101110010101;
            14'b10_100100110000: DATA = 12'b101110011000;
            14'b10_100100110001: DATA = 12'b101110011011;
            14'b10_100100110010: DATA = 12'b101110011101;
            14'b10_100100110011: DATA = 12'b101110100000;
            14'b10_100100110100: DATA = 12'b101110100011;
            14'b10_100100110101: DATA = 12'b101110100110;
            14'b10_100100110110: DATA = 12'b101110101001;
            14'b10_100100110111: DATA = 12'b101110101011;
            14'b10_100100111000: DATA = 12'b101110101110;
            14'b10_100100111001: DATA = 12'b101110110001;
            14'b10_100100111010: DATA = 12'b101110110100;
            14'b10_100100111011: DATA = 12'b101110110111;
            14'b10_100100111100: DATA = 12'b101110111001;
            14'b10_100100111101: DATA = 12'b101110111100;
            14'b10_100100111110: DATA = 12'b101110111111;
            14'b10_100100111111: DATA = 12'b101111000010;
            14'b10_100101000000: DATA = 12'b101111000100;
            14'b10_100101000001: DATA = 12'b101111000111;
            14'b10_100101000010: DATA = 12'b101111001010;
            14'b10_100101000011: DATA = 12'b101111001101;
            14'b10_100101000100: DATA = 12'b101111010000;
            14'b10_100101000101: DATA = 12'b101111010010;
            14'b10_100101000110: DATA = 12'b101111010101;
            14'b10_100101000111: DATA = 12'b101111011000;
            14'b10_100101001000: DATA = 12'b101111011011;
            14'b10_100101001001: DATA = 12'b101111011101;
            14'b10_100101001010: DATA = 12'b101111100000;
            14'b10_100101001011: DATA = 12'b101111100011;
            14'b10_100101001100: DATA = 12'b101111100110;
            14'b10_100101001101: DATA = 12'b101111101000;
            14'b10_100101001110: DATA = 12'b101111101011;
            14'b10_100101001111: DATA = 12'b101111101110;
            14'b10_100101010000: DATA = 12'b101111110000;
            14'b10_100101010001: DATA = 12'b101111110011;
            14'b10_100101010010: DATA = 12'b101111110110;
            14'b10_100101010011: DATA = 12'b101111111001;
            14'b10_100101010100: DATA = 12'b101111111011;
            14'b10_100101010101: DATA = 12'b101111111110;
            14'b10_100101010110: DATA = 12'b110000000001;
            14'b10_100101010111: DATA = 12'b110000000100;
            14'b10_100101011000: DATA = 12'b110000000110;
            14'b10_100101011001: DATA = 12'b110000001001;
            14'b10_100101011010: DATA = 12'b110000001100;
            14'b10_100101011011: DATA = 12'b110000001110;
            14'b10_100101011100: DATA = 12'b110000010001;
            14'b10_100101011101: DATA = 12'b110000010100;
            14'b10_100101011110: DATA = 12'b110000010110;
            14'b10_100101011111: DATA = 12'b110000011001;
            14'b10_100101100000: DATA = 12'b110000011100;
            14'b10_100101100001: DATA = 12'b110000011111;
            14'b10_100101100010: DATA = 12'b110000100001;
            14'b10_100101100011: DATA = 12'b110000100100;
            14'b10_100101100100: DATA = 12'b110000100111;
            14'b10_100101100101: DATA = 12'b110000101001;
            14'b10_100101100110: DATA = 12'b110000101100;
            14'b10_100101100111: DATA = 12'b110000101111;
            14'b10_100101101000: DATA = 12'b110000110001;
            14'b10_100101101001: DATA = 12'b110000110100;
            14'b10_100101101010: DATA = 12'b110000110111;
            14'b10_100101101011: DATA = 12'b110000111001;
            14'b10_100101101100: DATA = 12'b110000111100;
            14'b10_100101101101: DATA = 12'b110000111111;
            14'b10_100101101110: DATA = 12'b110001000001;
            14'b10_100101101111: DATA = 12'b110001000100;
            14'b10_100101110000: DATA = 12'b110001000111;
            14'b10_100101110001: DATA = 12'b110001001001;
            14'b10_100101110010: DATA = 12'b110001001100;
            14'b10_100101110011: DATA = 12'b110001001111;
            14'b10_100101110100: DATA = 12'b110001010001;
            14'b10_100101110101: DATA = 12'b110001010100;
            14'b10_100101110110: DATA = 12'b110001010111;
            14'b10_100101110111: DATA = 12'b110001011001;
            14'b10_100101111000: DATA = 12'b110001011100;
            14'b10_100101111001: DATA = 12'b110001011110;
            14'b10_100101111010: DATA = 12'b110001100001;
            14'b10_100101111011: DATA = 12'b110001100100;
            14'b10_100101111100: DATA = 12'b110001100110;
            14'b10_100101111101: DATA = 12'b110001101001;
            14'b10_100101111110: DATA = 12'b110001101100;
            14'b10_100101111111: DATA = 12'b110001101110;
            14'b10_100110000000: DATA = 12'b110001110001;
            14'b10_100110000001: DATA = 12'b110001110011;
            14'b10_100110000010: DATA = 12'b110001110110;
            14'b10_100110000011: DATA = 12'b110001111001;
            14'b10_100110000100: DATA = 12'b110001111011;
            14'b10_100110000101: DATA = 12'b110001111110;
            14'b10_100110000110: DATA = 12'b110010000000;
            14'b10_100110000111: DATA = 12'b110010000011;
            14'b10_100110001000: DATA = 12'b110010000110;
            14'b10_100110001001: DATA = 12'b110010001000;
            14'b10_100110001010: DATA = 12'b110010001011;
            14'b10_100110001011: DATA = 12'b110010001101;
            14'b10_100110001100: DATA = 12'b110010010000;
            14'b10_100110001101: DATA = 12'b110010010010;
            14'b10_100110001110: DATA = 12'b110010010101;
            14'b10_100110001111: DATA = 12'b110010011000;
            14'b10_100110010000: DATA = 12'b110010011010;
            14'b10_100110010001: DATA = 12'b110010011101;
            14'b10_100110010010: DATA = 12'b110010011111;
            14'b10_100110010011: DATA = 12'b110010100010;
            14'b10_100110010100: DATA = 12'b110010100100;
            14'b10_100110010101: DATA = 12'b110010100111;
            14'b10_100110010110: DATA = 12'b110010101010;
            14'b10_100110010111: DATA = 12'b110010101100;
            14'b10_100110011000: DATA = 12'b110010101111;
            14'b10_100110011001: DATA = 12'b110010110001;
            14'b10_100110011010: DATA = 12'b110010110100;
            14'b10_100110011011: DATA = 12'b110010110110;
            14'b10_100110011100: DATA = 12'b110010111001;
            14'b10_100110011101: DATA = 12'b110010111011;
            14'b10_100110011110: DATA = 12'b110010111110;
            14'b10_100110011111: DATA = 12'b110011000000;
            14'b10_100110100000: DATA = 12'b110011000011;
            14'b10_100110100001: DATA = 12'b110011000101;
            14'b10_100110100010: DATA = 12'b110011001000;
            14'b10_100110100011: DATA = 12'b110011001010;
            14'b10_100110100100: DATA = 12'b110011001101;
            14'b10_100110100101: DATA = 12'b110011001111;
            14'b10_100110100110: DATA = 12'b110011010010;
            14'b10_100110100111: DATA = 12'b110011010100;
            14'b10_100110101000: DATA = 12'b110011010111;
            14'b10_100110101001: DATA = 12'b110011011001;
            14'b10_100110101010: DATA = 12'b110011011100;
            14'b10_100110101011: DATA = 12'b110011011110;
            14'b10_100110101100: DATA = 12'b110011100001;
            14'b10_100110101101: DATA = 12'b110011100011;
            14'b10_100110101110: DATA = 12'b110011100110;
            14'b10_100110101111: DATA = 12'b110011101000;
            14'b10_100110110000: DATA = 12'b110011101011;
            14'b10_100110110001: DATA = 12'b110011101101;
            14'b10_100110110010: DATA = 12'b110011110000;
            14'b10_100110110011: DATA = 12'b110011110010;
            14'b10_100110110100: DATA = 12'b110011110101;
            14'b10_100110110101: DATA = 12'b110011110111;
            14'b10_100110110110: DATA = 12'b110011111010;
            14'b10_100110110111: DATA = 12'b110011111100;
            14'b10_100110111000: DATA = 12'b110011111111;
            14'b10_100110111001: DATA = 12'b110100000001;
            14'b10_100110111010: DATA = 12'b110100000011;
            14'b10_100110111011: DATA = 12'b110100000110;
            14'b10_100110111100: DATA = 12'b110100001000;
            14'b10_100110111101: DATA = 12'b110100001011;
            14'b10_100110111110: DATA = 12'b110100001101;
            14'b10_100110111111: DATA = 12'b110100010000;
            14'b10_100111000000: DATA = 12'b110100010010;
            14'b10_100111000001: DATA = 12'b110100010101;
            14'b10_100111000010: DATA = 12'b110100010111;
            14'b10_100111000011: DATA = 12'b110100011001;
            14'b10_100111000100: DATA = 12'b110100011100;
            14'b10_100111000101: DATA = 12'b110100011110;
            14'b10_100111000110: DATA = 12'b110100100001;
            14'b10_100111000111: DATA = 12'b110100100011;
            14'b10_100111001000: DATA = 12'b110100100101;
            14'b10_100111001001: DATA = 12'b110100101000;
            14'b10_100111001010: DATA = 12'b110100101010;
            14'b10_100111001011: DATA = 12'b110100101101;
            14'b10_100111001100: DATA = 12'b110100101111;
            14'b10_100111001101: DATA = 12'b110100110001;
            14'b10_100111001110: DATA = 12'b110100110100;
            14'b10_100111001111: DATA = 12'b110100110110;
            14'b10_100111010000: DATA = 12'b110100111001;
            14'b10_100111010001: DATA = 12'b110100111011;
            14'b10_100111010010: DATA = 12'b110100111101;
            14'b10_100111010011: DATA = 12'b110101000000;
            14'b10_100111010100: DATA = 12'b110101000010;
            14'b10_100111010101: DATA = 12'b110101000100;
            14'b10_100111010110: DATA = 12'b110101000111;
            14'b10_100111010111: DATA = 12'b110101001001;
            14'b10_100111011000: DATA = 12'b110101001011;
            14'b10_100111011001: DATA = 12'b110101001110;
            14'b10_100111011010: DATA = 12'b110101010000;
            14'b10_100111011011: DATA = 12'b110101010011;
            14'b10_100111011100: DATA = 12'b110101010101;
            14'b10_100111011101: DATA = 12'b110101010111;
            14'b10_100111011110: DATA = 12'b110101011010;
            14'b10_100111011111: DATA = 12'b110101011100;
            14'b10_100111100000: DATA = 12'b110101011110;
            14'b10_100111100001: DATA = 12'b110101100001;
            14'b10_100111100010: DATA = 12'b110101100011;
            14'b10_100111100011: DATA = 12'b110101100101;
            14'b10_100111100100: DATA = 12'b110101100111;
            14'b10_100111100101: DATA = 12'b110101101010;
            14'b10_100111100110: DATA = 12'b110101101100;
            14'b10_100111100111: DATA = 12'b110101101110;
            14'b10_100111101000: DATA = 12'b110101110001;
            14'b10_100111101001: DATA = 12'b110101110011;
            14'b10_100111101010: DATA = 12'b110101110101;
            14'b10_100111101011: DATA = 12'b110101111000;
            14'b10_100111101100: DATA = 12'b110101111010;
            14'b10_100111101101: DATA = 12'b110101111100;
            14'b10_100111101110: DATA = 12'b110101111110;
            14'b10_100111101111: DATA = 12'b110110000001;
            14'b10_100111110000: DATA = 12'b110110000011;
            14'b10_100111110001: DATA = 12'b110110000101;
            14'b10_100111110010: DATA = 12'b110110001000;
            14'b10_100111110011: DATA = 12'b110110001010;
            14'b10_100111110100: DATA = 12'b110110001100;
            14'b10_100111110101: DATA = 12'b110110001110;
            14'b10_100111110110: DATA = 12'b110110010001;
            14'b10_100111110111: DATA = 12'b110110010011;
            14'b10_100111111000: DATA = 12'b110110010101;
            14'b10_100111111001: DATA = 12'b110110010111;
            14'b10_100111111010: DATA = 12'b110110011010;
            14'b10_100111111011: DATA = 12'b110110011100;
            14'b10_100111111100: DATA = 12'b110110011110;
            14'b10_100111111101: DATA = 12'b110110100000;
            14'b10_100111111110: DATA = 12'b110110100011;
            14'b10_100111111111: DATA = 12'b110110100101;
            14'b10_101000000000: DATA = 12'b110110100111;
            14'b10_101000000001: DATA = 12'b110110101001;
            14'b10_101000000010: DATA = 12'b110110101011;
            14'b10_101000000011: DATA = 12'b110110101110;
            14'b10_101000000100: DATA = 12'b110110110000;
            14'b10_101000000101: DATA = 12'b110110110010;
            14'b10_101000000110: DATA = 12'b110110110100;
            14'b10_101000000111: DATA = 12'b110110110110;
            14'b10_101000001000: DATA = 12'b110110111001;
            14'b10_101000001001: DATA = 12'b110110111011;
            14'b10_101000001010: DATA = 12'b110110111101;
            14'b10_101000001011: DATA = 12'b110110111111;
            14'b10_101000001100: DATA = 12'b110111000001;
            14'b10_101000001101: DATA = 12'b110111000100;
            14'b10_101000001110: DATA = 12'b110111000110;
            14'b10_101000001111: DATA = 12'b110111001000;
            14'b10_101000010000: DATA = 12'b110111001010;
            14'b10_101000010001: DATA = 12'b110111001100;
            14'b10_101000010010: DATA = 12'b110111001110;
            14'b10_101000010011: DATA = 12'b110111010001;
            14'b10_101000010100: DATA = 12'b110111010011;
            14'b10_101000010101: DATA = 12'b110111010101;
            14'b10_101000010110: DATA = 12'b110111010111;
            14'b10_101000010111: DATA = 12'b110111011001;
            14'b10_101000011000: DATA = 12'b110111011011;
            14'b10_101000011001: DATA = 12'b110111011101;
            14'b10_101000011010: DATA = 12'b110111100000;
            14'b10_101000011011: DATA = 12'b110111100010;
            14'b10_101000011100: DATA = 12'b110111100100;
            14'b10_101000011101: DATA = 12'b110111100110;
            14'b10_101000011110: DATA = 12'b110111101000;
            14'b10_101000011111: DATA = 12'b110111101010;
            14'b10_101000100000: DATA = 12'b110111101100;
            14'b10_101000100001: DATA = 12'b110111101110;
            14'b10_101000100010: DATA = 12'b110111110000;
            14'b10_101000100011: DATA = 12'b110111110011;
            14'b10_101000100100: DATA = 12'b110111110101;
            14'b10_101000100101: DATA = 12'b110111110111;
            14'b10_101000100110: DATA = 12'b110111111001;
            14'b10_101000100111: DATA = 12'b110111111011;
            14'b10_101000101000: DATA = 12'b110111111101;
            14'b10_101000101001: DATA = 12'b110111111111;
            14'b10_101000101010: DATA = 12'b111000000001;
            14'b10_101000101011: DATA = 12'b111000000011;
            14'b10_101000101100: DATA = 12'b111000000101;
            14'b10_101000101101: DATA = 12'b111000000111;
            14'b10_101000101110: DATA = 12'b111000001001;
            14'b10_101000101111: DATA = 12'b111000001011;
            14'b10_101000110000: DATA = 12'b111000001110;
            14'b10_101000110001: DATA = 12'b111000010000;
            14'b10_101000110010: DATA = 12'b111000010010;
            14'b10_101000110011: DATA = 12'b111000010100;
            14'b10_101000110100: DATA = 12'b111000010110;
            14'b10_101000110101: DATA = 12'b111000011000;
            14'b10_101000110110: DATA = 12'b111000011010;
            14'b10_101000110111: DATA = 12'b111000011100;
            14'b10_101000111000: DATA = 12'b111000011110;
            14'b10_101000111001: DATA = 12'b111000100000;
            14'b10_101000111010: DATA = 12'b111000100010;
            14'b10_101000111011: DATA = 12'b111000100100;
            14'b10_101000111100: DATA = 12'b111000100110;
            14'b10_101000111101: DATA = 12'b111000101000;
            14'b10_101000111110: DATA = 12'b111000101010;
            14'b10_101000111111: DATA = 12'b111000101100;
            14'b10_101001000000: DATA = 12'b111000101110;
            14'b10_101001000001: DATA = 12'b111000110000;
            14'b10_101001000010: DATA = 12'b111000110010;
            14'b10_101001000011: DATA = 12'b111000110100;
            14'b10_101001000100: DATA = 12'b111000110110;
            14'b10_101001000101: DATA = 12'b111000111000;
            14'b10_101001000110: DATA = 12'b111000111010;
            14'b10_101001000111: DATA = 12'b111000111100;
            14'b10_101001001000: DATA = 12'b111000111110;
            14'b10_101001001001: DATA = 12'b111001000000;
            14'b10_101001001010: DATA = 12'b111001000010;
            14'b10_101001001011: DATA = 12'b111001000100;
            14'b10_101001001100: DATA = 12'b111001000101;
            14'b10_101001001101: DATA = 12'b111001000111;
            14'b10_101001001110: DATA = 12'b111001001001;
            14'b10_101001001111: DATA = 12'b111001001011;
            14'b10_101001010000: DATA = 12'b111001001101;
            14'b10_101001010001: DATA = 12'b111001001111;
            14'b10_101001010010: DATA = 12'b111001010001;
            14'b10_101001010011: DATA = 12'b111001010011;
            14'b10_101001010100: DATA = 12'b111001010101;
            14'b10_101001010101: DATA = 12'b111001010111;
            14'b10_101001010110: DATA = 12'b111001011001;
            14'b10_101001010111: DATA = 12'b111001011011;
            14'b10_101001011000: DATA = 12'b111001011101;
            14'b10_101001011001: DATA = 12'b111001011110;
            14'b10_101001011010: DATA = 12'b111001100000;
            14'b10_101001011011: DATA = 12'b111001100010;
            14'b10_101001011100: DATA = 12'b111001100100;
            14'b10_101001011101: DATA = 12'b111001100110;
            14'b10_101001011110: DATA = 12'b111001101000;
            14'b10_101001011111: DATA = 12'b111001101010;
            14'b10_101001100000: DATA = 12'b111001101100;
            14'b10_101001100001: DATA = 12'b111001101110;
            14'b10_101001100010: DATA = 12'b111001101111;
            14'b10_101001100011: DATA = 12'b111001110001;
            14'b10_101001100100: DATA = 12'b111001110011;
            14'b10_101001100101: DATA = 12'b111001110101;
            14'b10_101001100110: DATA = 12'b111001110111;
            14'b10_101001100111: DATA = 12'b111001111001;
            14'b10_101001101000: DATA = 12'b111001111011;
            14'b10_101001101001: DATA = 12'b111001111100;
            14'b10_101001101010: DATA = 12'b111001111110;
            14'b10_101001101011: DATA = 12'b111010000000;
            14'b10_101001101100: DATA = 12'b111010000010;
            14'b10_101001101101: DATA = 12'b111010000100;
            14'b10_101001101110: DATA = 12'b111010000101;
            14'b10_101001101111: DATA = 12'b111010000111;
            14'b10_101001110000: DATA = 12'b111010001001;
            14'b10_101001110001: DATA = 12'b111010001011;
            14'b10_101001110010: DATA = 12'b111010001101;
            14'b10_101001110011: DATA = 12'b111010001111;
            14'b10_101001110100: DATA = 12'b111010010000;
            14'b10_101001110101: DATA = 12'b111010010010;
            14'b10_101001110110: DATA = 12'b111010010100;
            14'b10_101001110111: DATA = 12'b111010010110;
            14'b10_101001111000: DATA = 12'b111010010111;
            14'b10_101001111001: DATA = 12'b111010011001;
            14'b10_101001111010: DATA = 12'b111010011011;
            14'b10_101001111011: DATA = 12'b111010011101;
            14'b10_101001111100: DATA = 12'b111010011111;
            14'b10_101001111101: DATA = 12'b111010100000;
            14'b10_101001111110: DATA = 12'b111010100010;
            14'b10_101001111111: DATA = 12'b111010100100;
            14'b10_101010000000: DATA = 12'b111010100110;
            14'b10_101010000001: DATA = 12'b111010100111;
            14'b10_101010000010: DATA = 12'b111010101001;
            14'b10_101010000011: DATA = 12'b111010101011;
            14'b10_101010000100: DATA = 12'b111010101100;
            14'b10_101010000101: DATA = 12'b111010101110;
            14'b10_101010000110: DATA = 12'b111010110000;
            14'b10_101010000111: DATA = 12'b111010110010;
            14'b10_101010001000: DATA = 12'b111010110011;
            14'b10_101010001001: DATA = 12'b111010110101;
            14'b10_101010001010: DATA = 12'b111010110111;
            14'b10_101010001011: DATA = 12'b111010111000;
            14'b10_101010001100: DATA = 12'b111010111010;
            14'b10_101010001101: DATA = 12'b111010111100;
            14'b10_101010001110: DATA = 12'b111010111110;
            14'b10_101010001111: DATA = 12'b111010111111;
            14'b10_101010010000: DATA = 12'b111011000001;
            14'b10_101010010001: DATA = 12'b111011000011;
            14'b10_101010010010: DATA = 12'b111011000100;
            14'b10_101010010011: DATA = 12'b111011000110;
            14'b10_101010010100: DATA = 12'b111011001000;
            14'b10_101010010101: DATA = 12'b111011001001;
            14'b10_101010010110: DATA = 12'b111011001011;
            14'b10_101010010111: DATA = 12'b111011001101;
            14'b10_101010011000: DATA = 12'b111011001110;
            14'b10_101010011001: DATA = 12'b111011010000;
            14'b10_101010011010: DATA = 12'b111011010010;
            14'b10_101010011011: DATA = 12'b111011010011;
            14'b10_101010011100: DATA = 12'b111011010101;
            14'b10_101010011101: DATA = 12'b111011010110;
            14'b10_101010011110: DATA = 12'b111011011000;
            14'b10_101010011111: DATA = 12'b111011011010;
            14'b10_101010100000: DATA = 12'b111011011011;
            14'b10_101010100001: DATA = 12'b111011011101;
            14'b10_101010100010: DATA = 12'b111011011110;
            14'b10_101010100011: DATA = 12'b111011100000;
            14'b10_101010100100: DATA = 12'b111011100010;
            14'b10_101010100101: DATA = 12'b111011100011;
            14'b10_101010100110: DATA = 12'b111011100101;
            14'b10_101010100111: DATA = 12'b111011100110;
            14'b10_101010101000: DATA = 12'b111011101000;
            14'b10_101010101001: DATA = 12'b111011101010;
            14'b10_101010101010: DATA = 12'b111011101011;
            14'b10_101010101011: DATA = 12'b111011101101;
            14'b10_101010101100: DATA = 12'b111011101110;
            14'b10_101010101101: DATA = 12'b111011110000;
            14'b10_101010101110: DATA = 12'b111011110001;
            14'b10_101010101111: DATA = 12'b111011110011;
            14'b10_101010110000: DATA = 12'b111011110101;
            14'b10_101010110001: DATA = 12'b111011110110;
            14'b10_101010110010: DATA = 12'b111011111000;
            14'b10_101010110011: DATA = 12'b111011111001;
            14'b10_101010110100: DATA = 12'b111011111011;
            14'b10_101010110101: DATA = 12'b111011111100;
            14'b10_101010110110: DATA = 12'b111011111110;
            14'b10_101010110111: DATA = 12'b111011111111;
            14'b10_101010111000: DATA = 12'b111100000001;
            14'b10_101010111001: DATA = 12'b111100000010;
            14'b10_101010111010: DATA = 12'b111100000100;
            14'b10_101010111011: DATA = 12'b111100000101;
            14'b10_101010111100: DATA = 12'b111100000111;
            14'b10_101010111101: DATA = 12'b111100001000;
            14'b10_101010111110: DATA = 12'b111100001010;
            14'b10_101010111111: DATA = 12'b111100001011;
            14'b10_101011000000: DATA = 12'b111100001101;
            14'b10_101011000001: DATA = 12'b111100001110;
            14'b10_101011000010: DATA = 12'b111100010000;
            14'b10_101011000011: DATA = 12'b111100010001;
            14'b10_101011000100: DATA = 12'b111100010011;
            14'b10_101011000101: DATA = 12'b111100010100;
            14'b10_101011000110: DATA = 12'b111100010110;
            14'b10_101011000111: DATA = 12'b111100010111;
            14'b10_101011001000: DATA = 12'b111100011000;
            14'b10_101011001001: DATA = 12'b111100011010;
            14'b10_101011001010: DATA = 12'b111100011011;
            14'b10_101011001011: DATA = 12'b111100011101;
            14'b10_101011001100: DATA = 12'b111100011110;
            14'b10_101011001101: DATA = 12'b111100100000;
            14'b10_101011001110: DATA = 12'b111100100001;
            14'b10_101011001111: DATA = 12'b111100100011;
            14'b10_101011010000: DATA = 12'b111100100100;
            14'b10_101011010001: DATA = 12'b111100100101;
            14'b10_101011010010: DATA = 12'b111100100111;
            14'b10_101011010011: DATA = 12'b111100101000;
            14'b10_101011010100: DATA = 12'b111100101010;
            14'b10_101011010101: DATA = 12'b111100101011;
            14'b10_101011010110: DATA = 12'b111100101100;
            14'b10_101011010111: DATA = 12'b111100101110;
            14'b10_101011011000: DATA = 12'b111100101111;
            14'b10_101011011001: DATA = 12'b111100110000;
            14'b10_101011011010: DATA = 12'b111100110010;
            14'b10_101011011011: DATA = 12'b111100110011;
            14'b10_101011011100: DATA = 12'b111100110101;
            14'b10_101011011101: DATA = 12'b111100110110;
            14'b10_101011011110: DATA = 12'b111100110111;
            14'b10_101011011111: DATA = 12'b111100111001;
            14'b10_101011100000: DATA = 12'b111100111010;
            14'b10_101011100001: DATA = 12'b111100111011;
            14'b10_101011100010: DATA = 12'b111100111101;
            14'b10_101011100011: DATA = 12'b111100111110;
            14'b10_101011100100: DATA = 12'b111100111111;
            14'b10_101011100101: DATA = 12'b111101000001;
            14'b10_101011100110: DATA = 12'b111101000010;
            14'b10_101011100111: DATA = 12'b111101000011;
            14'b10_101011101000: DATA = 12'b111101000101;
            14'b10_101011101001: DATA = 12'b111101000110;
            14'b10_101011101010: DATA = 12'b111101000111;
            14'b10_101011101011: DATA = 12'b111101001000;
            14'b10_101011101100: DATA = 12'b111101001010;
            14'b10_101011101101: DATA = 12'b111101001011;
            14'b10_101011101110: DATA = 12'b111101001100;
            14'b10_101011101111: DATA = 12'b111101001110;
            14'b10_101011110000: DATA = 12'b111101001111;
            14'b10_101011110001: DATA = 12'b111101010000;
            14'b10_101011110010: DATA = 12'b111101010001;
            14'b10_101011110011: DATA = 12'b111101010011;
            14'b10_101011110100: DATA = 12'b111101010100;
            14'b10_101011110101: DATA = 12'b111101010101;
            14'b10_101011110110: DATA = 12'b111101010110;
            14'b10_101011110111: DATA = 12'b111101011000;
            14'b10_101011111000: DATA = 12'b111101011001;
            14'b10_101011111001: DATA = 12'b111101011010;
            14'b10_101011111010: DATA = 12'b111101011011;
            14'b10_101011111011: DATA = 12'b111101011101;
            14'b10_101011111100: DATA = 12'b111101011110;
            14'b10_101011111101: DATA = 12'b111101011111;
            14'b10_101011111110: DATA = 12'b111101100000;
            14'b10_101011111111: DATA = 12'b111101100001;
            14'b10_101100000000: DATA = 12'b111101100011;
            14'b10_101100000001: DATA = 12'b111101100100;
            14'b10_101100000010: DATA = 12'b111101100101;
            14'b10_101100000011: DATA = 12'b111101100110;
            14'b10_101100000100: DATA = 12'b111101100111;
            14'b10_101100000101: DATA = 12'b111101101001;
            14'b10_101100000110: DATA = 12'b111101101010;
            14'b10_101100000111: DATA = 12'b111101101011;
            14'b10_101100001000: DATA = 12'b111101101100;
            14'b10_101100001001: DATA = 12'b111101101101;
            14'b10_101100001010: DATA = 12'b111101101110;
            14'b10_101100001011: DATA = 12'b111101110000;
            14'b10_101100001100: DATA = 12'b111101110001;
            14'b10_101100001101: DATA = 12'b111101110010;
            14'b10_101100001110: DATA = 12'b111101110011;
            14'b10_101100001111: DATA = 12'b111101110100;
            14'b10_101100010000: DATA = 12'b111101110101;
            14'b10_101100010001: DATA = 12'b111101110110;
            14'b10_101100010010: DATA = 12'b111101111000;
            14'b10_101100010011: DATA = 12'b111101111001;
            14'b10_101100010100: DATA = 12'b111101111010;
            14'b10_101100010101: DATA = 12'b111101111011;
            14'b10_101100010110: DATA = 12'b111101111100;
            14'b10_101100010111: DATA = 12'b111101111101;
            14'b10_101100011000: DATA = 12'b111101111110;
            14'b10_101100011001: DATA = 12'b111101111111;
            14'b10_101100011010: DATA = 12'b111110000000;
            14'b10_101100011011: DATA = 12'b111110000001;
            14'b10_101100011100: DATA = 12'b111110000011;
            14'b10_101100011101: DATA = 12'b111110000100;
            14'b10_101100011110: DATA = 12'b111110000101;
            14'b10_101100011111: DATA = 12'b111110000110;
            14'b10_101100100000: DATA = 12'b111110000111;
            14'b10_101100100001: DATA = 12'b111110001000;
            14'b10_101100100010: DATA = 12'b111110001001;
            14'b10_101100100011: DATA = 12'b111110001010;
            14'b10_101100100100: DATA = 12'b111110001011;
            14'b10_101100100101: DATA = 12'b111110001100;
            14'b10_101100100110: DATA = 12'b111110001101;
            14'b10_101100100111: DATA = 12'b111110001110;
            14'b10_101100101000: DATA = 12'b111110001111;
            14'b10_101100101001: DATA = 12'b111110010000;
            14'b10_101100101010: DATA = 12'b111110010001;
            14'b10_101100101011: DATA = 12'b111110010010;
            14'b10_101100101100: DATA = 12'b111110010011;
            14'b10_101100101101: DATA = 12'b111110010100;
            14'b10_101100101110: DATA = 12'b111110010101;
            14'b10_101100101111: DATA = 12'b111110010110;
            14'b10_101100110000: DATA = 12'b111110010111;
            14'b10_101100110001: DATA = 12'b111110011000;
            14'b10_101100110010: DATA = 12'b111110011001;
            14'b10_101100110011: DATA = 12'b111110011010;
            14'b10_101100110100: DATA = 12'b111110011011;
            14'b10_101100110101: DATA = 12'b111110011100;
            14'b10_101100110110: DATA = 12'b111110011101;
            14'b10_101100110111: DATA = 12'b111110011110;
            14'b10_101100111000: DATA = 12'b111110011111;
            14'b10_101100111001: DATA = 12'b111110100000;
            14'b10_101100111010: DATA = 12'b111110100001;
            14'b10_101100111011: DATA = 12'b111110100010;
            14'b10_101100111100: DATA = 12'b111110100011;
            14'b10_101100111101: DATA = 12'b111110100100;
            14'b10_101100111110: DATA = 12'b111110100101;
            14'b10_101100111111: DATA = 12'b111110100101;
            14'b10_101101000000: DATA = 12'b111110100110;
            14'b10_101101000001: DATA = 12'b111110100111;
            14'b10_101101000010: DATA = 12'b111110101000;
            14'b10_101101000011: DATA = 12'b111110101001;
            14'b10_101101000100: DATA = 12'b111110101010;
            14'b10_101101000101: DATA = 12'b111110101011;
            14'b10_101101000110: DATA = 12'b111110101100;
            14'b10_101101000111: DATA = 12'b111110101101;
            14'b10_101101001000: DATA = 12'b111110101110;
            14'b10_101101001001: DATA = 12'b111110101110;
            14'b10_101101001010: DATA = 12'b111110101111;
            14'b10_101101001011: DATA = 12'b111110110000;
            14'b10_101101001100: DATA = 12'b111110110001;
            14'b10_101101001101: DATA = 12'b111110110010;
            14'b10_101101001110: DATA = 12'b111110110011;
            14'b10_101101001111: DATA = 12'b111110110100;
            14'b10_101101010000: DATA = 12'b111110110100;
            14'b10_101101010001: DATA = 12'b111110110101;
            14'b10_101101010010: DATA = 12'b111110110110;
            14'b10_101101010011: DATA = 12'b111110110111;
            14'b10_101101010100: DATA = 12'b111110111000;
            14'b10_101101010101: DATA = 12'b111110111000;
            14'b10_101101010110: DATA = 12'b111110111001;
            14'b10_101101010111: DATA = 12'b111110111010;
            14'b10_101101011000: DATA = 12'b111110111011;
            14'b10_101101011001: DATA = 12'b111110111100;
            14'b10_101101011010: DATA = 12'b111110111100;
            14'b10_101101011011: DATA = 12'b111110111101;
            14'b10_101101011100: DATA = 12'b111110111110;
            14'b10_101101011101: DATA = 12'b111110111111;
            14'b10_101101011110: DATA = 12'b111111000000;
            14'b10_101101011111: DATA = 12'b111111000000;
            14'b10_101101100000: DATA = 12'b111111000001;
            14'b10_101101100001: DATA = 12'b111111000010;
            14'b10_101101100010: DATA = 12'b111111000011;
            14'b10_101101100011: DATA = 12'b111111000011;
            14'b10_101101100100: DATA = 12'b111111000100;
            14'b10_101101100101: DATA = 12'b111111000101;
            14'b10_101101100110: DATA = 12'b111111000110;
            14'b10_101101100111: DATA = 12'b111111000110;
            14'b10_101101101000: DATA = 12'b111111000111;
            14'b10_101101101001: DATA = 12'b111111001000;
            14'b10_101101101010: DATA = 12'b111111001001;
            14'b10_101101101011: DATA = 12'b111111001001;
            14'b10_101101101100: DATA = 12'b111111001010;
            14'b10_101101101101: DATA = 12'b111111001011;
            14'b10_101101101110: DATA = 12'b111111001011;
            14'b10_101101101111: DATA = 12'b111111001100;
            14'b10_101101110000: DATA = 12'b111111001101;
            14'b10_101101110001: DATA = 12'b111111001101;
            14'b10_101101110010: DATA = 12'b111111001110;
            14'b10_101101110011: DATA = 12'b111111001111;
            14'b10_101101110100: DATA = 12'b111111001111;
            14'b10_101101110101: DATA = 12'b111111010000;
            14'b10_101101110110: DATA = 12'b111111010001;
            14'b10_101101110111: DATA = 12'b111111010001;
            14'b10_101101111000: DATA = 12'b111111010010;
            14'b10_101101111001: DATA = 12'b111111010011;
            14'b10_101101111010: DATA = 12'b111111010011;
            14'b10_101101111011: DATA = 12'b111111010100;
            14'b10_101101111100: DATA = 12'b111111010101;
            14'b10_101101111101: DATA = 12'b111111010101;
            14'b10_101101111110: DATA = 12'b111111010110;
            14'b10_101101111111: DATA = 12'b111111010111;
            14'b10_101110000000: DATA = 12'b111111010111;
            14'b10_101110000001: DATA = 12'b111111011000;
            14'b10_101110000010: DATA = 12'b111111011000;
            14'b10_101110000011: DATA = 12'b111111011001;
            14'b10_101110000100: DATA = 12'b111111011010;
            14'b10_101110000101: DATA = 12'b111111011010;
            14'b10_101110000110: DATA = 12'b111111011011;
            14'b10_101110000111: DATA = 12'b111111011011;
            14'b10_101110001000: DATA = 12'b111111011100;
            14'b10_101110001001: DATA = 12'b111111011100;
            14'b10_101110001010: DATA = 12'b111111011101;
            14'b10_101110001011: DATA = 12'b111111011110;
            14'b10_101110001100: DATA = 12'b111111011110;
            14'b10_101110001101: DATA = 12'b111111011111;
            14'b10_101110001110: DATA = 12'b111111011111;
            14'b10_101110001111: DATA = 12'b111111100000;
            14'b10_101110010000: DATA = 12'b111111100000;
            14'b10_101110010001: DATA = 12'b111111100001;
            14'b10_101110010010: DATA = 12'b111111100001;
            14'b10_101110010011: DATA = 12'b111111100010;
            14'b10_101110010100: DATA = 12'b111111100010;
            14'b10_101110010101: DATA = 12'b111111100011;
            14'b10_101110010110: DATA = 12'b111111100011;
            14'b10_101110010111: DATA = 12'b111111100100;
            14'b10_101110011000: DATA = 12'b111111100101;
            14'b10_101110011001: DATA = 12'b111111100101;
            14'b10_101110011010: DATA = 12'b111111100101;
            14'b10_101110011011: DATA = 12'b111111100110;
            14'b10_101110011100: DATA = 12'b111111100110;
            14'b10_101110011101: DATA = 12'b111111100111;
            14'b10_101110011110: DATA = 12'b111111100111;
            14'b10_101110011111: DATA = 12'b111111101000;
            14'b10_101110100000: DATA = 12'b111111101000;
            14'b10_101110100001: DATA = 12'b111111101001;
            14'b10_101110100010: DATA = 12'b111111101001;
            14'b10_101110100011: DATA = 12'b111111101010;
            14'b10_101110100100: DATA = 12'b111111101010;
            14'b10_101110100101: DATA = 12'b111111101011;
            14'b10_101110100110: DATA = 12'b111111101011;
            14'b10_101110100111: DATA = 12'b111111101011;
            14'b10_101110101000: DATA = 12'b111111101100;
            14'b10_101110101001: DATA = 12'b111111101100;
            14'b10_101110101010: DATA = 12'b111111101101;
            14'b10_101110101011: DATA = 12'b111111101101;
            14'b10_101110101100: DATA = 12'b111111101110;
            14'b10_101110101101: DATA = 12'b111111101110;
            14'b10_101110101110: DATA = 12'b111111101110;
            14'b10_101110101111: DATA = 12'b111111101111;
            14'b10_101110110000: DATA = 12'b111111101111;
            14'b10_101110110001: DATA = 12'b111111101111;
            14'b10_101110110010: DATA = 12'b111111110000;
            14'b10_101110110011: DATA = 12'b111111110000;
            14'b10_101110110100: DATA = 12'b111111110001;
            14'b10_101110110101: DATA = 12'b111111110001;
            14'b10_101110110110: DATA = 12'b111111110001;
            14'b10_101110110111: DATA = 12'b111111110010;
            14'b10_101110111000: DATA = 12'b111111110010;
            14'b10_101110111001: DATA = 12'b111111110010;
            14'b10_101110111010: DATA = 12'b111111110011;
            14'b10_101110111011: DATA = 12'b111111110011;
            14'b10_101110111100: DATA = 12'b111111110011;
            14'b10_101110111101: DATA = 12'b111111110100;
            14'b10_101110111110: DATA = 12'b111111110100;
            14'b10_101110111111: DATA = 12'b111111110100;
            14'b10_101111000000: DATA = 12'b111111110101;
            14'b10_101111000001: DATA = 12'b111111110101;
            14'b10_101111000010: DATA = 12'b111111110101;
            14'b10_101111000011: DATA = 12'b111111110110;
            14'b10_101111000100: DATA = 12'b111111110110;
            14'b10_101111000101: DATA = 12'b111111110110;
            14'b10_101111000110: DATA = 12'b111111110110;
            14'b10_101111000111: DATA = 12'b111111110111;
            14'b10_101111001000: DATA = 12'b111111110111;
            14'b10_101111001001: DATA = 12'b111111110111;
            14'b10_101111001010: DATA = 12'b111111110111;
            14'b10_101111001011: DATA = 12'b111111111000;
            14'b10_101111001100: DATA = 12'b111111111000;
            14'b10_101111001101: DATA = 12'b111111111000;
            14'b10_101111001110: DATA = 12'b111111111000;
            14'b10_101111001111: DATA = 12'b111111111001;
            14'b10_101111010000: DATA = 12'b111111111001;
            14'b10_101111010001: DATA = 12'b111111111001;
            14'b10_101111010010: DATA = 12'b111111111001;
            14'b10_101111010011: DATA = 12'b111111111010;
            14'b10_101111010100: DATA = 12'b111111111010;
            14'b10_101111010101: DATA = 12'b111111111010;
            14'b10_101111010110: DATA = 12'b111111111010;
            14'b10_101111010111: DATA = 12'b111111111010;
            14'b10_101111011000: DATA = 12'b111111111011;
            14'b10_101111011001: DATA = 12'b111111111011;
            14'b10_101111011010: DATA = 12'b111111111011;
            14'b10_101111011011: DATA = 12'b111111111011;
            14'b10_101111011100: DATA = 12'b111111111011;
            14'b10_101111011101: DATA = 12'b111111111100;
            14'b10_101111011110: DATA = 12'b111111111100;
            14'b10_101111011111: DATA = 12'b111111111100;
            14'b10_101111100000: DATA = 12'b111111111100;
            14'b10_101111100001: DATA = 12'b111111111100;
            14'b10_101111100010: DATA = 12'b111111111100;
            14'b10_101111100011: DATA = 12'b111111111100;
            14'b10_101111100100: DATA = 12'b111111111101;
            14'b10_101111100101: DATA = 12'b111111111101;
            14'b10_101111100110: DATA = 12'b111111111101;
            14'b10_101111100111: DATA = 12'b111111111101;
            14'b10_101111101000: DATA = 12'b111111111101;
            14'b10_101111101001: DATA = 12'b111111111101;
            14'b10_101111101010: DATA = 12'b111111111101;
            14'b10_101111101011: DATA = 12'b111111111101;
            14'b10_101111101100: DATA = 12'b111111111110;
            14'b10_101111101101: DATA = 12'b111111111110;
            14'b10_101111101110: DATA = 12'b111111111110;
            14'b10_101111101111: DATA = 12'b111111111110;
            14'b10_101111110000: DATA = 12'b111111111110;
            14'b10_101111110001: DATA = 12'b111111111110;
            14'b10_101111110010: DATA = 12'b111111111110;
            14'b10_101111110011: DATA = 12'b111111111110;
            14'b10_101111110100: DATA = 12'b111111111110;
            14'b10_101111110101: DATA = 12'b111111111110;
            14'b10_101111110110: DATA = 12'b111111111110;
            14'b10_101111110111: DATA = 12'b111111111110;
            14'b10_101111111000: DATA = 12'b111111111110;
            14'b10_101111111001: DATA = 12'b111111111110;
            14'b10_101111111010: DATA = 12'b111111111110;
            14'b10_101111111011: DATA = 12'b111111111110;
            14'b10_101111111100: DATA = 12'b111111111110;
            14'b10_101111111101: DATA = 12'b111111111110;
            14'b10_101111111110: DATA = 12'b111111111110;
            14'b10_101111111111: DATA = 12'b111111111110;
            14'b10_110000000000: DATA = 12'b111111111111;
            14'b10_110000000001: DATA = 12'b111111111110;
            14'b10_110000000010: DATA = 12'b111111111110;
            14'b10_110000000011: DATA = 12'b111111111110;
            14'b10_110000000100: DATA = 12'b111111111110;
            14'b10_110000000101: DATA = 12'b111111111110;
            14'b10_110000000110: DATA = 12'b111111111110;
            14'b10_110000000111: DATA = 12'b111111111110;
            14'b10_110000001000: DATA = 12'b111111111110;
            14'b10_110000001001: DATA = 12'b111111111110;
            14'b10_110000001010: DATA = 12'b111111111110;
            14'b10_110000001011: DATA = 12'b111111111110;
            14'b10_110000001100: DATA = 12'b111111111110;
            14'b10_110000001101: DATA = 12'b111111111110;
            14'b10_110000001110: DATA = 12'b111111111110;
            14'b10_110000001111: DATA = 12'b111111111110;
            14'b10_110000010000: DATA = 12'b111111111110;
            14'b10_110000010001: DATA = 12'b111111111110;
            14'b10_110000010010: DATA = 12'b111111111110;
            14'b10_110000010011: DATA = 12'b111111111110;
            14'b10_110000010100: DATA = 12'b111111111110;
            14'b10_110000010101: DATA = 12'b111111111101;
            14'b10_110000010110: DATA = 12'b111111111101;
            14'b10_110000010111: DATA = 12'b111111111101;
            14'b10_110000011000: DATA = 12'b111111111101;
            14'b10_110000011001: DATA = 12'b111111111101;
            14'b10_110000011010: DATA = 12'b111111111101;
            14'b10_110000011011: DATA = 12'b111111111101;
            14'b10_110000011100: DATA = 12'b111111111101;
            14'b10_110000011101: DATA = 12'b111111111100;
            14'b10_110000011110: DATA = 12'b111111111100;
            14'b10_110000011111: DATA = 12'b111111111100;
            14'b10_110000100000: DATA = 12'b111111111100;
            14'b10_110000100001: DATA = 12'b111111111100;
            14'b10_110000100010: DATA = 12'b111111111100;
            14'b10_110000100011: DATA = 12'b111111111100;
            14'b10_110000100100: DATA = 12'b111111111011;
            14'b10_110000100101: DATA = 12'b111111111011;
            14'b10_110000100110: DATA = 12'b111111111011;
            14'b10_110000100111: DATA = 12'b111111111011;
            14'b10_110000101000: DATA = 12'b111111111011;
            14'b10_110000101001: DATA = 12'b111111111010;
            14'b10_110000101010: DATA = 12'b111111111010;
            14'b10_110000101011: DATA = 12'b111111111010;
            14'b10_110000101100: DATA = 12'b111111111010;
            14'b10_110000101101: DATA = 12'b111111111010;
            14'b10_110000101110: DATA = 12'b111111111001;
            14'b10_110000101111: DATA = 12'b111111111001;
            14'b10_110000110000: DATA = 12'b111111111001;
            14'b10_110000110001: DATA = 12'b111111111001;
            14'b10_110000110010: DATA = 12'b111111111000;
            14'b10_110000110011: DATA = 12'b111111111000;
            14'b10_110000110100: DATA = 12'b111111111000;
            14'b10_110000110101: DATA = 12'b111111111000;
            14'b10_110000110110: DATA = 12'b111111110111;
            14'b10_110000110111: DATA = 12'b111111110111;
            14'b10_110000111000: DATA = 12'b111111110111;
            14'b10_110000111001: DATA = 12'b111111110111;
            14'b10_110000111010: DATA = 12'b111111110110;
            14'b10_110000111011: DATA = 12'b111111110110;
            14'b10_110000111100: DATA = 12'b111111110110;
            14'b10_110000111101: DATA = 12'b111111110110;
            14'b10_110000111110: DATA = 12'b111111110101;
            14'b10_110000111111: DATA = 12'b111111110101;
            14'b10_110001000000: DATA = 12'b111111110101;
            14'b10_110001000001: DATA = 12'b111111110100;
            14'b10_110001000010: DATA = 12'b111111110100;
            14'b10_110001000011: DATA = 12'b111111110100;
            14'b10_110001000100: DATA = 12'b111111110011;
            14'b10_110001000101: DATA = 12'b111111110011;
            14'b10_110001000110: DATA = 12'b111111110011;
            14'b10_110001000111: DATA = 12'b111111110010;
            14'b10_110001001000: DATA = 12'b111111110010;
            14'b10_110001001001: DATA = 12'b111111110010;
            14'b10_110001001010: DATA = 12'b111111110001;
            14'b10_110001001011: DATA = 12'b111111110001;
            14'b10_110001001100: DATA = 12'b111111110001;
            14'b10_110001001101: DATA = 12'b111111110000;
            14'b10_110001001110: DATA = 12'b111111110000;
            14'b10_110001001111: DATA = 12'b111111101111;
            14'b10_110001010000: DATA = 12'b111111101111;
            14'b10_110001010001: DATA = 12'b111111101111;
            14'b10_110001010010: DATA = 12'b111111101110;
            14'b10_110001010011: DATA = 12'b111111101110;
            14'b10_110001010100: DATA = 12'b111111101110;
            14'b10_110001010101: DATA = 12'b111111101101;
            14'b10_110001010110: DATA = 12'b111111101101;
            14'b10_110001010111: DATA = 12'b111111101100;
            14'b10_110001011000: DATA = 12'b111111101100;
            14'b10_110001011001: DATA = 12'b111111101011;
            14'b10_110001011010: DATA = 12'b111111101011;
            14'b10_110001011011: DATA = 12'b111111101011;
            14'b10_110001011100: DATA = 12'b111111101010;
            14'b10_110001011101: DATA = 12'b111111101010;
            14'b10_110001011110: DATA = 12'b111111101001;
            14'b10_110001011111: DATA = 12'b111111101001;
            14'b10_110001100000: DATA = 12'b111111101000;
            14'b10_110001100001: DATA = 12'b111111101000;
            14'b10_110001100010: DATA = 12'b111111100111;
            14'b10_110001100011: DATA = 12'b111111100111;
            14'b10_110001100100: DATA = 12'b111111100110;
            14'b10_110001100101: DATA = 12'b111111100110;
            14'b10_110001100110: DATA = 12'b111111100101;
            14'b10_110001100111: DATA = 12'b111111100101;
            14'b10_110001101000: DATA = 12'b111111100101;
            14'b10_110001101001: DATA = 12'b111111100100;
            14'b10_110001101010: DATA = 12'b111111100011;
            14'b10_110001101011: DATA = 12'b111111100011;
            14'b10_110001101100: DATA = 12'b111111100010;
            14'b10_110001101101: DATA = 12'b111111100010;
            14'b10_110001101110: DATA = 12'b111111100001;
            14'b10_110001101111: DATA = 12'b111111100001;
            14'b10_110001110000: DATA = 12'b111111100000;
            14'b10_110001110001: DATA = 12'b111111100000;
            14'b10_110001110010: DATA = 12'b111111011111;
            14'b10_110001110011: DATA = 12'b111111011111;
            14'b10_110001110100: DATA = 12'b111111011110;
            14'b10_110001110101: DATA = 12'b111111011110;
            14'b10_110001110110: DATA = 12'b111111011101;
            14'b10_110001110111: DATA = 12'b111111011100;
            14'b10_110001111000: DATA = 12'b111111011100;
            14'b10_110001111001: DATA = 12'b111111011011;
            14'b10_110001111010: DATA = 12'b111111011011;
            14'b10_110001111011: DATA = 12'b111111011010;
            14'b10_110001111100: DATA = 12'b111111011010;
            14'b10_110001111101: DATA = 12'b111111011001;
            14'b10_110001111110: DATA = 12'b111111011000;
            14'b10_110001111111: DATA = 12'b111111011000;
            14'b10_110010000000: DATA = 12'b111111010111;
            14'b10_110010000001: DATA = 12'b111111010111;
            14'b10_110010000010: DATA = 12'b111111010110;
            14'b10_110010000011: DATA = 12'b111111010101;
            14'b10_110010000100: DATA = 12'b111111010101;
            14'b10_110010000101: DATA = 12'b111111010100;
            14'b10_110010000110: DATA = 12'b111111010011;
            14'b10_110010000111: DATA = 12'b111111010011;
            14'b10_110010001000: DATA = 12'b111111010010;
            14'b10_110010001001: DATA = 12'b111111010001;
            14'b10_110010001010: DATA = 12'b111111010001;
            14'b10_110010001011: DATA = 12'b111111010000;
            14'b10_110010001100: DATA = 12'b111111001111;
            14'b10_110010001101: DATA = 12'b111111001111;
            14'b10_110010001110: DATA = 12'b111111001110;
            14'b10_110010001111: DATA = 12'b111111001101;
            14'b10_110010010000: DATA = 12'b111111001101;
            14'b10_110010010001: DATA = 12'b111111001100;
            14'b10_110010010010: DATA = 12'b111111001011;
            14'b10_110010010011: DATA = 12'b111111001011;
            14'b10_110010010100: DATA = 12'b111111001010;
            14'b10_110010010101: DATA = 12'b111111001001;
            14'b10_110010010110: DATA = 12'b111111001001;
            14'b10_110010010111: DATA = 12'b111111001000;
            14'b10_110010011000: DATA = 12'b111111000111;
            14'b10_110010011001: DATA = 12'b111111000110;
            14'b10_110010011010: DATA = 12'b111111000110;
            14'b10_110010011011: DATA = 12'b111111000101;
            14'b10_110010011100: DATA = 12'b111111000100;
            14'b10_110010011101: DATA = 12'b111111000011;
            14'b10_110010011110: DATA = 12'b111111000011;
            14'b10_110010011111: DATA = 12'b111111000010;
            14'b10_110010100000: DATA = 12'b111111000001;
            14'b10_110010100001: DATA = 12'b111111000000;
            14'b10_110010100010: DATA = 12'b111111000000;
            14'b10_110010100011: DATA = 12'b111110111111;
            14'b10_110010100100: DATA = 12'b111110111110;
            14'b10_110010100101: DATA = 12'b111110111101;
            14'b10_110010100110: DATA = 12'b111110111100;
            14'b10_110010100111: DATA = 12'b111110111100;
            14'b10_110010101000: DATA = 12'b111110111011;
            14'b10_110010101001: DATA = 12'b111110111010;
            14'b10_110010101010: DATA = 12'b111110111001;
            14'b10_110010101011: DATA = 12'b111110111000;
            14'b10_110010101100: DATA = 12'b111110111000;
            14'b10_110010101101: DATA = 12'b111110110111;
            14'b10_110010101110: DATA = 12'b111110110110;
            14'b10_110010101111: DATA = 12'b111110110101;
            14'b10_110010110000: DATA = 12'b111110110100;
            14'b10_110010110001: DATA = 12'b111110110100;
            14'b10_110010110010: DATA = 12'b111110110011;
            14'b10_110010110011: DATA = 12'b111110110010;
            14'b10_110010110100: DATA = 12'b111110110001;
            14'b10_110010110101: DATA = 12'b111110110000;
            14'b10_110010110110: DATA = 12'b111110101111;
            14'b10_110010110111: DATA = 12'b111110101110;
            14'b10_110010111000: DATA = 12'b111110101110;
            14'b10_110010111001: DATA = 12'b111110101101;
            14'b10_110010111010: DATA = 12'b111110101100;
            14'b10_110010111011: DATA = 12'b111110101011;
            14'b10_110010111100: DATA = 12'b111110101010;
            14'b10_110010111101: DATA = 12'b111110101001;
            14'b10_110010111110: DATA = 12'b111110101000;
            14'b10_110010111111: DATA = 12'b111110100111;
            14'b10_110011000000: DATA = 12'b111110100110;
            14'b10_110011000001: DATA = 12'b111110100101;
            14'b10_110011000010: DATA = 12'b111110100101;
            14'b10_110011000011: DATA = 12'b111110100100;
            14'b10_110011000100: DATA = 12'b111110100011;
            14'b10_110011000101: DATA = 12'b111110100010;
            14'b10_110011000110: DATA = 12'b111110100001;
            14'b10_110011000111: DATA = 12'b111110100000;
            14'b10_110011001000: DATA = 12'b111110011111;
            14'b10_110011001001: DATA = 12'b111110011110;
            14'b10_110011001010: DATA = 12'b111110011101;
            14'b10_110011001011: DATA = 12'b111110011100;
            14'b10_110011001100: DATA = 12'b111110011011;
            14'b10_110011001101: DATA = 12'b111110011010;
            14'b10_110011001110: DATA = 12'b111110011001;
            14'b10_110011001111: DATA = 12'b111110011000;
            14'b10_110011010000: DATA = 12'b111110010111;
            14'b10_110011010001: DATA = 12'b111110010110;
            14'b10_110011010010: DATA = 12'b111110010101;
            14'b10_110011010011: DATA = 12'b111110010100;
            14'b10_110011010100: DATA = 12'b111110010011;
            14'b10_110011010101: DATA = 12'b111110010010;
            14'b10_110011010110: DATA = 12'b111110010001;
            14'b10_110011010111: DATA = 12'b111110010000;
            14'b10_110011011000: DATA = 12'b111110001111;
            14'b10_110011011001: DATA = 12'b111110001110;
            14'b10_110011011010: DATA = 12'b111110001101;
            14'b10_110011011011: DATA = 12'b111110001100;
            14'b10_110011011100: DATA = 12'b111110001011;
            14'b10_110011011101: DATA = 12'b111110001010;
            14'b10_110011011110: DATA = 12'b111110001001;
            14'b10_110011011111: DATA = 12'b111110001000;
            14'b10_110011100000: DATA = 12'b111110000111;
            14'b10_110011100001: DATA = 12'b111110000110;
            14'b10_110011100010: DATA = 12'b111110000101;
            14'b10_110011100011: DATA = 12'b111110000100;
            14'b10_110011100100: DATA = 12'b111110000011;
            14'b10_110011100101: DATA = 12'b111110000001;
            14'b10_110011100110: DATA = 12'b111110000000;
            14'b10_110011100111: DATA = 12'b111101111111;
            14'b10_110011101000: DATA = 12'b111101111110;
            14'b10_110011101001: DATA = 12'b111101111101;
            14'b10_110011101010: DATA = 12'b111101111100;
            14'b10_110011101011: DATA = 12'b111101111011;
            14'b10_110011101100: DATA = 12'b111101111010;
            14'b10_110011101101: DATA = 12'b111101111001;
            14'b10_110011101110: DATA = 12'b111101111000;
            14'b10_110011101111: DATA = 12'b111101110110;
            14'b10_110011110000: DATA = 12'b111101110101;
            14'b10_110011110001: DATA = 12'b111101110100;
            14'b10_110011110010: DATA = 12'b111101110011;
            14'b10_110011110011: DATA = 12'b111101110010;
            14'b10_110011110100: DATA = 12'b111101110001;
            14'b10_110011110101: DATA = 12'b111101110000;
            14'b10_110011110110: DATA = 12'b111101101110;
            14'b10_110011110111: DATA = 12'b111101101101;
            14'b10_110011111000: DATA = 12'b111101101100;
            14'b10_110011111001: DATA = 12'b111101101011;
            14'b10_110011111010: DATA = 12'b111101101010;
            14'b10_110011111011: DATA = 12'b111101101001;
            14'b10_110011111100: DATA = 12'b111101100111;
            14'b10_110011111101: DATA = 12'b111101100110;
            14'b10_110011111110: DATA = 12'b111101100101;
            14'b10_110011111111: DATA = 12'b111101100100;
            14'b10_110100000000: DATA = 12'b111101100011;
            14'b10_110100000001: DATA = 12'b111101100001;
            14'b10_110100000010: DATA = 12'b111101100000;
            14'b10_110100000011: DATA = 12'b111101011111;
            14'b10_110100000100: DATA = 12'b111101011110;
            14'b10_110100000101: DATA = 12'b111101011101;
            14'b10_110100000110: DATA = 12'b111101011011;
            14'b10_110100000111: DATA = 12'b111101011010;
            14'b10_110100001000: DATA = 12'b111101011001;
            14'b10_110100001001: DATA = 12'b111101011000;
            14'b10_110100001010: DATA = 12'b111101010110;
            14'b10_110100001011: DATA = 12'b111101010101;
            14'b10_110100001100: DATA = 12'b111101010100;
            14'b10_110100001101: DATA = 12'b111101010011;
            14'b10_110100001110: DATA = 12'b111101010001;
            14'b10_110100001111: DATA = 12'b111101010000;
            14'b10_110100010000: DATA = 12'b111101001111;
            14'b10_110100010001: DATA = 12'b111101001110;
            14'b10_110100010010: DATA = 12'b111101001100;
            14'b10_110100010011: DATA = 12'b111101001011;
            14'b10_110100010100: DATA = 12'b111101001010;
            14'b10_110100010101: DATA = 12'b111101001000;
            14'b10_110100010110: DATA = 12'b111101000111;
            14'b10_110100010111: DATA = 12'b111101000110;
            14'b10_110100011000: DATA = 12'b111101000101;
            14'b10_110100011001: DATA = 12'b111101000011;
            14'b10_110100011010: DATA = 12'b111101000010;
            14'b10_110100011011: DATA = 12'b111101000001;
            14'b10_110100011100: DATA = 12'b111100111111;
            14'b10_110100011101: DATA = 12'b111100111110;
            14'b10_110100011110: DATA = 12'b111100111101;
            14'b10_110100011111: DATA = 12'b111100111011;
            14'b10_110100100000: DATA = 12'b111100111010;
            14'b10_110100100001: DATA = 12'b111100111001;
            14'b10_110100100010: DATA = 12'b111100110111;
            14'b10_110100100011: DATA = 12'b111100110110;
            14'b10_110100100100: DATA = 12'b111100110101;
            14'b10_110100100101: DATA = 12'b111100110011;
            14'b10_110100100110: DATA = 12'b111100110010;
            14'b10_110100100111: DATA = 12'b111100110000;
            14'b10_110100101000: DATA = 12'b111100101111;
            14'b10_110100101001: DATA = 12'b111100101110;
            14'b10_110100101010: DATA = 12'b111100101100;
            14'b10_110100101011: DATA = 12'b111100101011;
            14'b10_110100101100: DATA = 12'b111100101010;
            14'b10_110100101101: DATA = 12'b111100101000;
            14'b10_110100101110: DATA = 12'b111100100111;
            14'b10_110100101111: DATA = 12'b111100100101;
            14'b10_110100110000: DATA = 12'b111100100100;
            14'b10_110100110001: DATA = 12'b111100100011;
            14'b10_110100110010: DATA = 12'b111100100001;
            14'b10_110100110011: DATA = 12'b111100100000;
            14'b10_110100110100: DATA = 12'b111100011110;
            14'b10_110100110101: DATA = 12'b111100011101;
            14'b10_110100110110: DATA = 12'b111100011011;
            14'b10_110100110111: DATA = 12'b111100011010;
            14'b10_110100111000: DATA = 12'b111100011000;
            14'b10_110100111001: DATA = 12'b111100010111;
            14'b10_110100111010: DATA = 12'b111100010110;
            14'b10_110100111011: DATA = 12'b111100010100;
            14'b10_110100111100: DATA = 12'b111100010011;
            14'b10_110100111101: DATA = 12'b111100010001;
            14'b10_110100111110: DATA = 12'b111100010000;
            14'b10_110100111111: DATA = 12'b111100001110;
            14'b10_110101000000: DATA = 12'b111100001101;
            14'b10_110101000001: DATA = 12'b111100001011;
            14'b10_110101000010: DATA = 12'b111100001010;
            14'b10_110101000011: DATA = 12'b111100001000;
            14'b10_110101000100: DATA = 12'b111100000111;
            14'b10_110101000101: DATA = 12'b111100000101;
            14'b10_110101000110: DATA = 12'b111100000100;
            14'b10_110101000111: DATA = 12'b111100000010;
            14'b10_110101001000: DATA = 12'b111100000001;
            14'b10_110101001001: DATA = 12'b111011111111;
            14'b10_110101001010: DATA = 12'b111011111110;
            14'b10_110101001011: DATA = 12'b111011111100;
            14'b10_110101001100: DATA = 12'b111011111011;
            14'b10_110101001101: DATA = 12'b111011111001;
            14'b10_110101001110: DATA = 12'b111011111000;
            14'b10_110101001111: DATA = 12'b111011110110;
            14'b10_110101010000: DATA = 12'b111011110101;
            14'b10_110101010001: DATA = 12'b111011110011;
            14'b10_110101010010: DATA = 12'b111011110001;
            14'b10_110101010011: DATA = 12'b111011110000;
            14'b10_110101010100: DATA = 12'b111011101110;
            14'b10_110101010101: DATA = 12'b111011101101;
            14'b10_110101010110: DATA = 12'b111011101011;
            14'b10_110101010111: DATA = 12'b111011101010;
            14'b10_110101011000: DATA = 12'b111011101000;
            14'b10_110101011001: DATA = 12'b111011100110;
            14'b10_110101011010: DATA = 12'b111011100101;
            14'b10_110101011011: DATA = 12'b111011100011;
            14'b10_110101011100: DATA = 12'b111011100010;
            14'b10_110101011101: DATA = 12'b111011100000;
            14'b10_110101011110: DATA = 12'b111011011110;
            14'b10_110101011111: DATA = 12'b111011011101;
            14'b10_110101100000: DATA = 12'b111011011011;
            14'b10_110101100001: DATA = 12'b111011011010;
            14'b10_110101100010: DATA = 12'b111011011000;
            14'b10_110101100011: DATA = 12'b111011010110;
            14'b10_110101100100: DATA = 12'b111011010101;
            14'b10_110101100101: DATA = 12'b111011010011;
            14'b10_110101100110: DATA = 12'b111011010010;
            14'b10_110101100111: DATA = 12'b111011010000;
            14'b10_110101101000: DATA = 12'b111011001110;
            14'b10_110101101001: DATA = 12'b111011001101;
            14'b10_110101101010: DATA = 12'b111011001011;
            14'b10_110101101011: DATA = 12'b111011001001;
            14'b10_110101101100: DATA = 12'b111011001000;
            14'b10_110101101101: DATA = 12'b111011000110;
            14'b10_110101101110: DATA = 12'b111011000100;
            14'b10_110101101111: DATA = 12'b111011000011;
            14'b10_110101110000: DATA = 12'b111011000001;
            14'b10_110101110001: DATA = 12'b111010111111;
            14'b10_110101110010: DATA = 12'b111010111110;
            14'b10_110101110011: DATA = 12'b111010111100;
            14'b10_110101110100: DATA = 12'b111010111010;
            14'b10_110101110101: DATA = 12'b111010111000;
            14'b10_110101110110: DATA = 12'b111010110111;
            14'b10_110101110111: DATA = 12'b111010110101;
            14'b10_110101111000: DATA = 12'b111010110011;
            14'b10_110101111001: DATA = 12'b111010110010;
            14'b10_110101111010: DATA = 12'b111010110000;
            14'b10_110101111011: DATA = 12'b111010101110;
            14'b10_110101111100: DATA = 12'b111010101100;
            14'b10_110101111101: DATA = 12'b111010101011;
            14'b10_110101111110: DATA = 12'b111010101001;
            14'b10_110101111111: DATA = 12'b111010100111;
            14'b10_110110000000: DATA = 12'b111010100110;
            14'b10_110110000001: DATA = 12'b111010100100;
            14'b10_110110000010: DATA = 12'b111010100010;
            14'b10_110110000011: DATA = 12'b111010100000;
            14'b10_110110000100: DATA = 12'b111010011111;
            14'b10_110110000101: DATA = 12'b111010011101;
            14'b10_110110000110: DATA = 12'b111010011011;
            14'b10_110110000111: DATA = 12'b111010011001;
            14'b10_110110001000: DATA = 12'b111010010111;
            14'b10_110110001001: DATA = 12'b111010010110;
            14'b10_110110001010: DATA = 12'b111010010100;
            14'b10_110110001011: DATA = 12'b111010010010;
            14'b10_110110001100: DATA = 12'b111010010000;
            14'b10_110110001101: DATA = 12'b111010001111;
            14'b10_110110001110: DATA = 12'b111010001101;
            14'b10_110110001111: DATA = 12'b111010001011;
            14'b10_110110010000: DATA = 12'b111010001001;
            14'b10_110110010001: DATA = 12'b111010000111;
            14'b10_110110010010: DATA = 12'b111010000101;
            14'b10_110110010011: DATA = 12'b111010000100;
            14'b10_110110010100: DATA = 12'b111010000010;
            14'b10_110110010101: DATA = 12'b111010000000;
            14'b10_110110010110: DATA = 12'b111001111110;
            14'b10_110110010111: DATA = 12'b111001111100;
            14'b10_110110011000: DATA = 12'b111001111011;
            14'b10_110110011001: DATA = 12'b111001111001;
            14'b10_110110011010: DATA = 12'b111001110111;
            14'b10_110110011011: DATA = 12'b111001110101;
            14'b10_110110011100: DATA = 12'b111001110011;
            14'b10_110110011101: DATA = 12'b111001110001;
            14'b10_110110011110: DATA = 12'b111001101111;
            14'b10_110110011111: DATA = 12'b111001101110;
            14'b10_110110100000: DATA = 12'b111001101100;
            14'b10_110110100001: DATA = 12'b111001101010;
            14'b10_110110100010: DATA = 12'b111001101000;
            14'b10_110110100011: DATA = 12'b111001100110;
            14'b10_110110100100: DATA = 12'b111001100100;
            14'b10_110110100101: DATA = 12'b111001100010;
            14'b10_110110100110: DATA = 12'b111001100000;
            14'b10_110110100111: DATA = 12'b111001011110;
            14'b10_110110101000: DATA = 12'b111001011101;
            14'b10_110110101001: DATA = 12'b111001011011;
            14'b10_110110101010: DATA = 12'b111001011001;
            14'b10_110110101011: DATA = 12'b111001010111;
            14'b10_110110101100: DATA = 12'b111001010101;
            14'b10_110110101101: DATA = 12'b111001010011;
            14'b10_110110101110: DATA = 12'b111001010001;
            14'b10_110110101111: DATA = 12'b111001001111;
            14'b10_110110110000: DATA = 12'b111001001101;
            14'b10_110110110001: DATA = 12'b111001001011;
            14'b10_110110110010: DATA = 12'b111001001001;
            14'b10_110110110011: DATA = 12'b111001000111;
            14'b10_110110110100: DATA = 12'b111001000101;
            14'b10_110110110101: DATA = 12'b111001000100;
            14'b10_110110110110: DATA = 12'b111001000010;
            14'b10_110110110111: DATA = 12'b111001000000;
            14'b10_110110111000: DATA = 12'b111000111110;
            14'b10_110110111001: DATA = 12'b111000111100;
            14'b10_110110111010: DATA = 12'b111000111010;
            14'b10_110110111011: DATA = 12'b111000111000;
            14'b10_110110111100: DATA = 12'b111000110110;
            14'b10_110110111101: DATA = 12'b111000110100;
            14'b10_110110111110: DATA = 12'b111000110010;
            14'b10_110110111111: DATA = 12'b111000110000;
            14'b10_110111000000: DATA = 12'b111000101110;
            14'b10_110111000001: DATA = 12'b111000101100;
            14'b10_110111000010: DATA = 12'b111000101010;
            14'b10_110111000011: DATA = 12'b111000101000;
            14'b10_110111000100: DATA = 12'b111000100110;
            14'b10_110111000101: DATA = 12'b111000100100;
            14'b10_110111000110: DATA = 12'b111000100010;
            14'b10_110111000111: DATA = 12'b111000100000;
            14'b10_110111001000: DATA = 12'b111000011110;
            14'b10_110111001001: DATA = 12'b111000011100;
            14'b10_110111001010: DATA = 12'b111000011010;
            14'b10_110111001011: DATA = 12'b111000011000;
            14'b10_110111001100: DATA = 12'b111000010110;
            14'b10_110111001101: DATA = 12'b111000010100;
            14'b10_110111001110: DATA = 12'b111000010010;
            14'b10_110111001111: DATA = 12'b111000010000;
            14'b10_110111010000: DATA = 12'b111000001110;
            14'b10_110111010001: DATA = 12'b111000001011;
            14'b10_110111010010: DATA = 12'b111000001001;
            14'b10_110111010011: DATA = 12'b111000000111;
            14'b10_110111010100: DATA = 12'b111000000101;
            14'b10_110111010101: DATA = 12'b111000000011;
            14'b10_110111010110: DATA = 12'b111000000001;
            14'b10_110111010111: DATA = 12'b110111111111;
            14'b10_110111011000: DATA = 12'b110111111101;
            14'b10_110111011001: DATA = 12'b110111111011;
            14'b10_110111011010: DATA = 12'b110111111001;
            14'b10_110111011011: DATA = 12'b110111110111;
            14'b10_110111011100: DATA = 12'b110111110101;
            14'b10_110111011101: DATA = 12'b110111110011;
            14'b10_110111011110: DATA = 12'b110111110000;
            14'b10_110111011111: DATA = 12'b110111101110;
            14'b10_110111100000: DATA = 12'b110111101100;
            14'b10_110111100001: DATA = 12'b110111101010;
            14'b10_110111100010: DATA = 12'b110111101000;
            14'b10_110111100011: DATA = 12'b110111100110;
            14'b10_110111100100: DATA = 12'b110111100100;
            14'b10_110111100101: DATA = 12'b110111100010;
            14'b10_110111100110: DATA = 12'b110111100000;
            14'b10_110111100111: DATA = 12'b110111011101;
            14'b10_110111101000: DATA = 12'b110111011011;
            14'b10_110111101001: DATA = 12'b110111011001;
            14'b10_110111101010: DATA = 12'b110111010111;
            14'b10_110111101011: DATA = 12'b110111010101;
            14'b10_110111101100: DATA = 12'b110111010011;
            14'b10_110111101101: DATA = 12'b110111010001;
            14'b10_110111101110: DATA = 12'b110111001110;
            14'b10_110111101111: DATA = 12'b110111001100;
            14'b10_110111110000: DATA = 12'b110111001010;
            14'b10_110111110001: DATA = 12'b110111001000;
            14'b10_110111110010: DATA = 12'b110111000110;
            14'b10_110111110011: DATA = 12'b110111000100;
            14'b10_110111110100: DATA = 12'b110111000001;
            14'b10_110111110101: DATA = 12'b110110111111;
            14'b10_110111110110: DATA = 12'b110110111101;
            14'b10_110111110111: DATA = 12'b110110111011;
            14'b10_110111111000: DATA = 12'b110110111001;
            14'b10_110111111001: DATA = 12'b110110110110;
            14'b10_110111111010: DATA = 12'b110110110100;
            14'b10_110111111011: DATA = 12'b110110110010;
            14'b10_110111111100: DATA = 12'b110110110000;
            14'b10_110111111101: DATA = 12'b110110101110;
            14'b10_110111111110: DATA = 12'b110110101011;
            14'b10_110111111111: DATA = 12'b110110101001;
            14'b10_111000000000: DATA = 12'b110110100111;
            14'b10_111000000001: DATA = 12'b110110100101;
            14'b10_111000000010: DATA = 12'b110110100011;
            14'b10_111000000011: DATA = 12'b110110100000;
            14'b10_111000000100: DATA = 12'b110110011110;
            14'b10_111000000101: DATA = 12'b110110011100;
            14'b10_111000000110: DATA = 12'b110110011010;
            14'b10_111000000111: DATA = 12'b110110010111;
            14'b10_111000001000: DATA = 12'b110110010101;
            14'b10_111000001001: DATA = 12'b110110010011;
            14'b10_111000001010: DATA = 12'b110110010001;
            14'b10_111000001011: DATA = 12'b110110001110;
            14'b10_111000001100: DATA = 12'b110110001100;
            14'b10_111000001101: DATA = 12'b110110001010;
            14'b10_111000001110: DATA = 12'b110110001000;
            14'b10_111000001111: DATA = 12'b110110000101;
            14'b10_111000010000: DATA = 12'b110110000011;
            14'b10_111000010001: DATA = 12'b110110000001;
            14'b10_111000010010: DATA = 12'b110101111110;
            14'b10_111000010011: DATA = 12'b110101111100;
            14'b10_111000010100: DATA = 12'b110101111010;
            14'b10_111000010101: DATA = 12'b110101111000;
            14'b10_111000010110: DATA = 12'b110101110101;
            14'b10_111000010111: DATA = 12'b110101110011;
            14'b10_111000011000: DATA = 12'b110101110001;
            14'b10_111000011001: DATA = 12'b110101101110;
            14'b10_111000011010: DATA = 12'b110101101100;
            14'b10_111000011011: DATA = 12'b110101101010;
            14'b10_111000011100: DATA = 12'b110101100111;
            14'b10_111000011101: DATA = 12'b110101100101;
            14'b10_111000011110: DATA = 12'b110101100011;
            14'b10_111000011111: DATA = 12'b110101100001;
            14'b10_111000100000: DATA = 12'b110101011110;
            14'b10_111000100001: DATA = 12'b110101011100;
            14'b10_111000100010: DATA = 12'b110101011010;
            14'b10_111000100011: DATA = 12'b110101010111;
            14'b10_111000100100: DATA = 12'b110101010101;
            14'b10_111000100101: DATA = 12'b110101010011;
            14'b10_111000100110: DATA = 12'b110101010000;
            14'b10_111000100111: DATA = 12'b110101001110;
            14'b10_111000101000: DATA = 12'b110101001011;
            14'b10_111000101001: DATA = 12'b110101001001;
            14'b10_111000101010: DATA = 12'b110101000111;
            14'b10_111000101011: DATA = 12'b110101000100;
            14'b10_111000101100: DATA = 12'b110101000010;
            14'b10_111000101101: DATA = 12'b110101000000;
            14'b10_111000101110: DATA = 12'b110100111101;
            14'b10_111000101111: DATA = 12'b110100111011;
            14'b10_111000110000: DATA = 12'b110100111001;
            14'b10_111000110001: DATA = 12'b110100110110;
            14'b10_111000110010: DATA = 12'b110100110100;
            14'b10_111000110011: DATA = 12'b110100110001;
            14'b10_111000110100: DATA = 12'b110100101111;
            14'b10_111000110101: DATA = 12'b110100101101;
            14'b10_111000110110: DATA = 12'b110100101010;
            14'b10_111000110111: DATA = 12'b110100101000;
            14'b10_111000111000: DATA = 12'b110100100101;
            14'b10_111000111001: DATA = 12'b110100100011;
            14'b10_111000111010: DATA = 12'b110100100001;
            14'b10_111000111011: DATA = 12'b110100011110;
            14'b10_111000111100: DATA = 12'b110100011100;
            14'b10_111000111101: DATA = 12'b110100011001;
            14'b10_111000111110: DATA = 12'b110100010111;
            14'b10_111000111111: DATA = 12'b110100010101;
            14'b10_111001000000: DATA = 12'b110100010010;
            14'b10_111001000001: DATA = 12'b110100010000;
            14'b10_111001000010: DATA = 12'b110100001101;
            14'b10_111001000011: DATA = 12'b110100001011;
            14'b10_111001000100: DATA = 12'b110100001000;
            14'b10_111001000101: DATA = 12'b110100000110;
            14'b10_111001000110: DATA = 12'b110100000011;
            14'b10_111001000111: DATA = 12'b110100000001;
            14'b10_111001001000: DATA = 12'b110011111111;
            14'b10_111001001001: DATA = 12'b110011111100;
            14'b10_111001001010: DATA = 12'b110011111010;
            14'b10_111001001011: DATA = 12'b110011110111;
            14'b10_111001001100: DATA = 12'b110011110101;
            14'b10_111001001101: DATA = 12'b110011110010;
            14'b10_111001001110: DATA = 12'b110011110000;
            14'b10_111001001111: DATA = 12'b110011101101;
            14'b10_111001010000: DATA = 12'b110011101011;
            14'b10_111001010001: DATA = 12'b110011101000;
            14'b10_111001010010: DATA = 12'b110011100110;
            14'b10_111001010011: DATA = 12'b110011100011;
            14'b10_111001010100: DATA = 12'b110011100001;
            14'b10_111001010101: DATA = 12'b110011011110;
            14'b10_111001010110: DATA = 12'b110011011100;
            14'b10_111001010111: DATA = 12'b110011011001;
            14'b10_111001011000: DATA = 12'b110011010111;
            14'b10_111001011001: DATA = 12'b110011010100;
            14'b10_111001011010: DATA = 12'b110011010010;
            14'b10_111001011011: DATA = 12'b110011001111;
            14'b10_111001011100: DATA = 12'b110011001101;
            14'b10_111001011101: DATA = 12'b110011001010;
            14'b10_111001011110: DATA = 12'b110011001000;
            14'b10_111001011111: DATA = 12'b110011000101;
            14'b10_111001100000: DATA = 12'b110011000011;
            14'b10_111001100001: DATA = 12'b110011000000;
            14'b10_111001100010: DATA = 12'b110010111110;
            14'b10_111001100011: DATA = 12'b110010111011;
            14'b10_111001100100: DATA = 12'b110010111001;
            14'b10_111001100101: DATA = 12'b110010110110;
            14'b10_111001100110: DATA = 12'b110010110100;
            14'b10_111001100111: DATA = 12'b110010110001;
            14'b10_111001101000: DATA = 12'b110010101111;
            14'b10_111001101001: DATA = 12'b110010101100;
            14'b10_111001101010: DATA = 12'b110010101010;
            14'b10_111001101011: DATA = 12'b110010100111;
            14'b10_111001101100: DATA = 12'b110010100100;
            14'b10_111001101101: DATA = 12'b110010100010;
            14'b10_111001101110: DATA = 12'b110010011111;
            14'b10_111001101111: DATA = 12'b110010011101;
            14'b10_111001110000: DATA = 12'b110010011010;
            14'b10_111001110001: DATA = 12'b110010011000;
            14'b10_111001110010: DATA = 12'b110010010101;
            14'b10_111001110011: DATA = 12'b110010010010;
            14'b10_111001110100: DATA = 12'b110010010000;
            14'b10_111001110101: DATA = 12'b110010001101;
            14'b10_111001110110: DATA = 12'b110010001011;
            14'b10_111001110111: DATA = 12'b110010001000;
            14'b10_111001111000: DATA = 12'b110010000110;
            14'b10_111001111001: DATA = 12'b110010000011;
            14'b10_111001111010: DATA = 12'b110010000000;
            14'b10_111001111011: DATA = 12'b110001111110;
            14'b10_111001111100: DATA = 12'b110001111011;
            14'b10_111001111101: DATA = 12'b110001111001;
            14'b10_111001111110: DATA = 12'b110001110110;
            14'b10_111001111111: DATA = 12'b110001110011;
            14'b10_111010000000: DATA = 12'b110001110001;
            14'b10_111010000001: DATA = 12'b110001101110;
            14'b10_111010000010: DATA = 12'b110001101100;
            14'b10_111010000011: DATA = 12'b110001101001;
            14'b10_111010000100: DATA = 12'b110001100110;
            14'b10_111010000101: DATA = 12'b110001100100;
            14'b10_111010000110: DATA = 12'b110001100001;
            14'b10_111010000111: DATA = 12'b110001011110;
            14'b10_111010001000: DATA = 12'b110001011100;
            14'b10_111010001001: DATA = 12'b110001011001;
            14'b10_111010001010: DATA = 12'b110001010111;
            14'b10_111010001011: DATA = 12'b110001010100;
            14'b10_111010001100: DATA = 12'b110001010001;
            14'b10_111010001101: DATA = 12'b110001001111;
            14'b10_111010001110: DATA = 12'b110001001100;
            14'b10_111010001111: DATA = 12'b110001001001;
            14'b10_111010010000: DATA = 12'b110001000111;
            14'b10_111010010001: DATA = 12'b110001000100;
            14'b10_111010010010: DATA = 12'b110001000001;
            14'b10_111010010011: DATA = 12'b110000111111;
            14'b10_111010010100: DATA = 12'b110000111100;
            14'b10_111010010101: DATA = 12'b110000111001;
            14'b10_111010010110: DATA = 12'b110000110111;
            14'b10_111010010111: DATA = 12'b110000110100;
            14'b10_111010011000: DATA = 12'b110000110001;
            14'b10_111010011001: DATA = 12'b110000101111;
            14'b10_111010011010: DATA = 12'b110000101100;
            14'b10_111010011011: DATA = 12'b110000101001;
            14'b10_111010011100: DATA = 12'b110000100111;
            14'b10_111010011101: DATA = 12'b110000100100;
            14'b10_111010011110: DATA = 12'b110000100001;
            14'b10_111010011111: DATA = 12'b110000011111;
            14'b10_111010100000: DATA = 12'b110000011100;
            14'b10_111010100001: DATA = 12'b110000011001;
            14'b10_111010100010: DATA = 12'b110000010110;
            14'b10_111010100011: DATA = 12'b110000010100;
            14'b10_111010100100: DATA = 12'b110000010001;
            14'b10_111010100101: DATA = 12'b110000001110;
            14'b10_111010100110: DATA = 12'b110000001100;
            14'b10_111010100111: DATA = 12'b110000001001;
            14'b10_111010101000: DATA = 12'b110000000110;
            14'b10_111010101001: DATA = 12'b110000000100;
            14'b10_111010101010: DATA = 12'b110000000001;
            14'b10_111010101011: DATA = 12'b101111111110;
            14'b10_111010101100: DATA = 12'b101111111011;
            14'b10_111010101101: DATA = 12'b101111111001;
            14'b10_111010101110: DATA = 12'b101111110110;
            14'b10_111010101111: DATA = 12'b101111110011;
            14'b10_111010110000: DATA = 12'b101111110000;
            14'b10_111010110001: DATA = 12'b101111101110;
            14'b10_111010110010: DATA = 12'b101111101011;
            14'b10_111010110011: DATA = 12'b101111101000;
            14'b10_111010110100: DATA = 12'b101111100110;
            14'b10_111010110101: DATA = 12'b101111100011;
            14'b10_111010110110: DATA = 12'b101111100000;
            14'b10_111010110111: DATA = 12'b101111011101;
            14'b10_111010111000: DATA = 12'b101111011011;
            14'b10_111010111001: DATA = 12'b101111011000;
            14'b10_111010111010: DATA = 12'b101111010101;
            14'b10_111010111011: DATA = 12'b101111010010;
            14'b10_111010111100: DATA = 12'b101111010000;
            14'b10_111010111101: DATA = 12'b101111001101;
            14'b10_111010111110: DATA = 12'b101111001010;
            14'b10_111010111111: DATA = 12'b101111000111;
            14'b10_111011000000: DATA = 12'b101111000100;
            14'b10_111011000001: DATA = 12'b101111000010;
            14'b10_111011000010: DATA = 12'b101110111111;
            14'b10_111011000011: DATA = 12'b101110111100;
            14'b10_111011000100: DATA = 12'b101110111001;
            14'b10_111011000101: DATA = 12'b101110110111;
            14'b10_111011000110: DATA = 12'b101110110100;
            14'b10_111011000111: DATA = 12'b101110110001;
            14'b10_111011001000: DATA = 12'b101110101110;
            14'b10_111011001001: DATA = 12'b101110101011;
            14'b10_111011001010: DATA = 12'b101110101001;
            14'b10_111011001011: DATA = 12'b101110100110;
            14'b10_111011001100: DATA = 12'b101110100011;
            14'b10_111011001101: DATA = 12'b101110100000;
            14'b10_111011001110: DATA = 12'b101110011101;
            14'b10_111011001111: DATA = 12'b101110011011;
            14'b10_111011010000: DATA = 12'b101110011000;
            14'b10_111011010001: DATA = 12'b101110010101;
            14'b10_111011010010: DATA = 12'b101110010010;
            14'b10_111011010011: DATA = 12'b101110001111;
            14'b10_111011010100: DATA = 12'b101110001101;
            14'b10_111011010101: DATA = 12'b101110001010;
            14'b10_111011010110: DATA = 12'b101110000111;
            14'b10_111011010111: DATA = 12'b101110000100;
            14'b10_111011011000: DATA = 12'b101110000001;
            14'b10_111011011001: DATA = 12'b101101111111;
            14'b10_111011011010: DATA = 12'b101101111100;
            14'b10_111011011011: DATA = 12'b101101111001;
            14'b10_111011011100: DATA = 12'b101101110110;
            14'b10_111011011101: DATA = 12'b101101110011;
            14'b10_111011011110: DATA = 12'b101101110000;
            14'b10_111011011111: DATA = 12'b101101101110;
            14'b10_111011100000: DATA = 12'b101101101011;
            14'b10_111011100001: DATA = 12'b101101101000;
            14'b10_111011100010: DATA = 12'b101101100101;
            14'b10_111011100011: DATA = 12'b101101100010;
            14'b10_111011100100: DATA = 12'b101101011111;
            14'b10_111011100101: DATA = 12'b101101011100;
            14'b10_111011100110: DATA = 12'b101101011010;
            14'b10_111011100111: DATA = 12'b101101010111;
            14'b10_111011101000: DATA = 12'b101101010100;
            14'b10_111011101001: DATA = 12'b101101010001;
            14'b10_111011101010: DATA = 12'b101101001110;
            14'b10_111011101011: DATA = 12'b101101001011;
            14'b10_111011101100: DATA = 12'b101101001000;
            14'b10_111011101101: DATA = 12'b101101000110;
            14'b10_111011101110: DATA = 12'b101101000011;
            14'b10_111011101111: DATA = 12'b101101000000;
            14'b10_111011110000: DATA = 12'b101100111101;
            14'b10_111011110001: DATA = 12'b101100111010;
            14'b10_111011110010: DATA = 12'b101100110111;
            14'b10_111011110011: DATA = 12'b101100110100;
            14'b10_111011110100: DATA = 12'b101100110010;
            14'b10_111011110101: DATA = 12'b101100101111;
            14'b10_111011110110: DATA = 12'b101100101100;
            14'b10_111011110111: DATA = 12'b101100101001;
            14'b10_111011111000: DATA = 12'b101100100110;
            14'b10_111011111001: DATA = 12'b101100100011;
            14'b10_111011111010: DATA = 12'b101100100000;
            14'b10_111011111011: DATA = 12'b101100011101;
            14'b10_111011111100: DATA = 12'b101100011010;
            14'b10_111011111101: DATA = 12'b101100011000;
            14'b10_111011111110: DATA = 12'b101100010101;
            14'b10_111011111111: DATA = 12'b101100010010;
            14'b10_111100000000: DATA = 12'b101100001111;
            14'b10_111100000001: DATA = 12'b101100001100;
            14'b10_111100000010: DATA = 12'b101100001001;
            14'b10_111100000011: DATA = 12'b101100000110;
            14'b10_111100000100: DATA = 12'b101100000011;
            14'b10_111100000101: DATA = 12'b101100000000;
            14'b10_111100000110: DATA = 12'b101011111101;
            14'b10_111100000111: DATA = 12'b101011111011;
            14'b10_111100001000: DATA = 12'b101011111000;
            14'b10_111100001001: DATA = 12'b101011110101;
            14'b10_111100001010: DATA = 12'b101011110010;
            14'b10_111100001011: DATA = 12'b101011101111;
            14'b10_111100001100: DATA = 12'b101011101100;
            14'b10_111100001101: DATA = 12'b101011101001;
            14'b10_111100001110: DATA = 12'b101011100110;
            14'b10_111100001111: DATA = 12'b101011100011;
            14'b10_111100010000: DATA = 12'b101011100000;
            14'b10_111100010001: DATA = 12'b101011011101;
            14'b10_111100010010: DATA = 12'b101011011010;
            14'b10_111100010011: DATA = 12'b101011010111;
            14'b10_111100010100: DATA = 12'b101011010100;
            14'b10_111100010101: DATA = 12'b101011010010;
            14'b10_111100010110: DATA = 12'b101011001111;
            14'b10_111100010111: DATA = 12'b101011001100;
            14'b10_111100011000: DATA = 12'b101011001001;
            14'b10_111100011001: DATA = 12'b101011000110;
            14'b10_111100011010: DATA = 12'b101011000011;
            14'b10_111100011011: DATA = 12'b101011000000;
            14'b10_111100011100: DATA = 12'b101010111101;
            14'b10_111100011101: DATA = 12'b101010111010;
            14'b10_111100011110: DATA = 12'b101010110111;
            14'b10_111100011111: DATA = 12'b101010110100;
            14'b10_111100100000: DATA = 12'b101010110001;
            14'b10_111100100001: DATA = 12'b101010101110;
            14'b10_111100100010: DATA = 12'b101010101011;
            14'b10_111100100011: DATA = 12'b101010101000;
            14'b10_111100100100: DATA = 12'b101010100101;
            14'b10_111100100101: DATA = 12'b101010100010;
            14'b10_111100100110: DATA = 12'b101010011111;
            14'b10_111100100111: DATA = 12'b101010011100;
            14'b10_111100101000: DATA = 12'b101010011001;
            14'b10_111100101001: DATA = 12'b101010010110;
            14'b10_111100101010: DATA = 12'b101010010011;
            14'b10_111100101011: DATA = 12'b101010010000;
            14'b10_111100101100: DATA = 12'b101010001110;
            14'b10_111100101101: DATA = 12'b101010001011;
            14'b10_111100101110: DATA = 12'b101010001000;
            14'b10_111100101111: DATA = 12'b101010000101;
            14'b10_111100110000: DATA = 12'b101010000010;
            14'b10_111100110001: DATA = 12'b101001111111;
            14'b10_111100110010: DATA = 12'b101001111100;
            14'b10_111100110011: DATA = 12'b101001111001;
            14'b10_111100110100: DATA = 12'b101001110110;
            14'b10_111100110101: DATA = 12'b101001110011;
            14'b10_111100110110: DATA = 12'b101001110000;
            14'b10_111100110111: DATA = 12'b101001101101;
            14'b10_111100111000: DATA = 12'b101001101010;
            14'b10_111100111001: DATA = 12'b101001100111;
            14'b10_111100111010: DATA = 12'b101001100100;
            14'b10_111100111011: DATA = 12'b101001100001;
            14'b10_111100111100: DATA = 12'b101001011110;
            14'b10_111100111101: DATA = 12'b101001011011;
            14'b10_111100111110: DATA = 12'b101001011000;
            14'b10_111100111111: DATA = 12'b101001010101;
            14'b10_111101000000: DATA = 12'b101001010010;
            14'b10_111101000001: DATA = 12'b101001001111;
            14'b10_111101000010: DATA = 12'b101001001100;
            14'b10_111101000011: DATA = 12'b101001001001;
            14'b10_111101000100: DATA = 12'b101001000110;
            14'b10_111101000101: DATA = 12'b101001000011;
            14'b10_111101000110: DATA = 12'b101001000000;
            14'b10_111101000111: DATA = 12'b101000111101;
            14'b10_111101001000: DATA = 12'b101000111010;
            14'b10_111101001001: DATA = 12'b101000110111;
            14'b10_111101001010: DATA = 12'b101000110100;
            14'b10_111101001011: DATA = 12'b101000110001;
            14'b10_111101001100: DATA = 12'b101000101110;
            14'b10_111101001101: DATA = 12'b101000101011;
            14'b10_111101001110: DATA = 12'b101000101000;
            14'b10_111101001111: DATA = 12'b101000100100;
            14'b10_111101010000: DATA = 12'b101000100001;
            14'b10_111101010001: DATA = 12'b101000011110;
            14'b10_111101010010: DATA = 12'b101000011011;
            14'b10_111101010011: DATA = 12'b101000011000;
            14'b10_111101010100: DATA = 12'b101000010101;
            14'b10_111101010101: DATA = 12'b101000010010;
            14'b10_111101010110: DATA = 12'b101000001111;
            14'b10_111101010111: DATA = 12'b101000001100;
            14'b10_111101011000: DATA = 12'b101000001001;
            14'b10_111101011001: DATA = 12'b101000000110;
            14'b10_111101011010: DATA = 12'b101000000011;
            14'b10_111101011011: DATA = 12'b101000000000;
            14'b10_111101011100: DATA = 12'b100111111101;
            14'b10_111101011101: DATA = 12'b100111111010;
            14'b10_111101011110: DATA = 12'b100111110111;
            14'b10_111101011111: DATA = 12'b100111110100;
            14'b10_111101100000: DATA = 12'b100111110001;
            14'b10_111101100001: DATA = 12'b100111101110;
            14'b10_111101100010: DATA = 12'b100111101011;
            14'b10_111101100011: DATA = 12'b100111101000;
            14'b10_111101100100: DATA = 12'b100111100101;
            14'b10_111101100101: DATA = 12'b100111100010;
            14'b10_111101100110: DATA = 12'b100111011111;
            14'b10_111101100111: DATA = 12'b100111011100;
            14'b10_111101101000: DATA = 12'b100111011000;
            14'b10_111101101001: DATA = 12'b100111010101;
            14'b10_111101101010: DATA = 12'b100111010010;
            14'b10_111101101011: DATA = 12'b100111001111;
            14'b10_111101101100: DATA = 12'b100111001100;
            14'b10_111101101101: DATA = 12'b100111001001;
            14'b10_111101101110: DATA = 12'b100111000110;
            14'b10_111101101111: DATA = 12'b100111000011;
            14'b10_111101110000: DATA = 12'b100111000000;
            14'b10_111101110001: DATA = 12'b100110111101;
            14'b10_111101110010: DATA = 12'b100110111010;
            14'b10_111101110011: DATA = 12'b100110110111;
            14'b10_111101110100: DATA = 12'b100110110100;
            14'b10_111101110101: DATA = 12'b100110110001;
            14'b10_111101110110: DATA = 12'b100110101110;
            14'b10_111101110111: DATA = 12'b100110101011;
            14'b10_111101111000: DATA = 12'b100110100111;
            14'b10_111101111001: DATA = 12'b100110100100;
            14'b10_111101111010: DATA = 12'b100110100001;
            14'b10_111101111011: DATA = 12'b100110011110;
            14'b10_111101111100: DATA = 12'b100110011011;
            14'b10_111101111101: DATA = 12'b100110011000;
            14'b10_111101111110: DATA = 12'b100110010101;
            14'b10_111101111111: DATA = 12'b100110010010;
            14'b10_111110000000: DATA = 12'b100110001111;
            14'b10_111110000001: DATA = 12'b100110001100;
            14'b10_111110000010: DATA = 12'b100110001001;
            14'b10_111110000011: DATA = 12'b100110000110;
            14'b10_111110000100: DATA = 12'b100110000011;
            14'b10_111110000101: DATA = 12'b100101111111;
            14'b10_111110000110: DATA = 12'b100101111100;
            14'b10_111110000111: DATA = 12'b100101111001;
            14'b10_111110001000: DATA = 12'b100101110110;
            14'b10_111110001001: DATA = 12'b100101110011;
            14'b10_111110001010: DATA = 12'b100101110000;
            14'b10_111110001011: DATA = 12'b100101101101;
            14'b10_111110001100: DATA = 12'b100101101010;
            14'b10_111110001101: DATA = 12'b100101100111;
            14'b10_111110001110: DATA = 12'b100101100100;
            14'b10_111110001111: DATA = 12'b100101100001;
            14'b10_111110010000: DATA = 12'b100101011101;
            14'b10_111110010001: DATA = 12'b100101011010;
            14'b10_111110010010: DATA = 12'b100101010111;
            14'b10_111110010011: DATA = 12'b100101010100;
            14'b10_111110010100: DATA = 12'b100101010001;
            14'b10_111110010101: DATA = 12'b100101001110;
            14'b10_111110010110: DATA = 12'b100101001011;
            14'b10_111110010111: DATA = 12'b100101001000;
            14'b10_111110011000: DATA = 12'b100101000101;
            14'b10_111110011001: DATA = 12'b100101000010;
            14'b10_111110011010: DATA = 12'b100100111110;
            14'b10_111110011011: DATA = 12'b100100111011;
            14'b10_111110011100: DATA = 12'b100100111000;
            14'b10_111110011101: DATA = 12'b100100110101;
            14'b10_111110011110: DATA = 12'b100100110010;
            14'b10_111110011111: DATA = 12'b100100101111;
            14'b10_111110100000: DATA = 12'b100100101100;
            14'b10_111110100001: DATA = 12'b100100101001;
            14'b10_111110100010: DATA = 12'b100100100110;
            14'b10_111110100011: DATA = 12'b100100100011;
            14'b10_111110100100: DATA = 12'b100100011111;
            14'b10_111110100101: DATA = 12'b100100011100;
            14'b10_111110100110: DATA = 12'b100100011001;
            14'b10_111110100111: DATA = 12'b100100010110;
            14'b10_111110101000: DATA = 12'b100100010011;
            14'b10_111110101001: DATA = 12'b100100010000;
            14'b10_111110101010: DATA = 12'b100100001101;
            14'b10_111110101011: DATA = 12'b100100001010;
            14'b10_111110101100: DATA = 12'b100100000111;
            14'b10_111110101101: DATA = 12'b100100000011;
            14'b10_111110101110: DATA = 12'b100100000000;
            14'b10_111110101111: DATA = 12'b100011111101;
            14'b10_111110110000: DATA = 12'b100011111010;
            14'b10_111110110001: DATA = 12'b100011110111;
            14'b10_111110110010: DATA = 12'b100011110100;
            14'b10_111110110011: DATA = 12'b100011110001;
            14'b10_111110110100: DATA = 12'b100011101110;
            14'b10_111110110101: DATA = 12'b100011101010;
            14'b10_111110110110: DATA = 12'b100011100111;
            14'b10_111110110111: DATA = 12'b100011100100;
            14'b10_111110111000: DATA = 12'b100011100001;
            14'b10_111110111001: DATA = 12'b100011011110;
            14'b10_111110111010: DATA = 12'b100011011011;
            14'b10_111110111011: DATA = 12'b100011011000;
            14'b10_111110111100: DATA = 12'b100011010101;
            14'b10_111110111101: DATA = 12'b100011010010;
            14'b10_111110111110: DATA = 12'b100011001110;
            14'b10_111110111111: DATA = 12'b100011001011;
            14'b10_111111000000: DATA = 12'b100011001000;
            14'b10_111111000001: DATA = 12'b100011000101;
            14'b10_111111000010: DATA = 12'b100011000010;
            14'b10_111111000011: DATA = 12'b100010111111;
            14'b10_111111000100: DATA = 12'b100010111100;
            14'b10_111111000101: DATA = 12'b100010111001;
            14'b10_111111000110: DATA = 12'b100010110101;
            14'b10_111111000111: DATA = 12'b100010110010;
            14'b10_111111001000: DATA = 12'b100010101111;
            14'b10_111111001001: DATA = 12'b100010101100;
            14'b10_111111001010: DATA = 12'b100010101001;
            14'b10_111111001011: DATA = 12'b100010100110;
            14'b10_111111001100: DATA = 12'b100010100011;
            14'b10_111111001101: DATA = 12'b100010011111;
            14'b10_111111001110: DATA = 12'b100010011100;
            14'b10_111111001111: DATA = 12'b100010011001;
            14'b10_111111010000: DATA = 12'b100010010110;
            14'b10_111111010001: DATA = 12'b100010010011;
            14'b10_111111010010: DATA = 12'b100010010000;
            14'b10_111111010011: DATA = 12'b100010001101;
            14'b10_111111010100: DATA = 12'b100010001010;
            14'b10_111111010101: DATA = 12'b100010000110;
            14'b10_111111010110: DATA = 12'b100010000011;
            14'b10_111111010111: DATA = 12'b100010000000;
            14'b10_111111011000: DATA = 12'b100001111101;
            14'b10_111111011001: DATA = 12'b100001111010;
            14'b10_111111011010: DATA = 12'b100001110111;
            14'b10_111111011011: DATA = 12'b100001110100;
            14'b10_111111011100: DATA = 12'b100001110000;
            14'b10_111111011101: DATA = 12'b100001101101;
            14'b10_111111011110: DATA = 12'b100001101010;
            14'b10_111111011111: DATA = 12'b100001100111;
            14'b10_111111100000: DATA = 12'b100001100100;
            14'b10_111111100001: DATA = 12'b100001100001;
            14'b10_111111100010: DATA = 12'b100001011110;
            14'b10_111111100011: DATA = 12'b100001011011;
            14'b10_111111100100: DATA = 12'b100001010111;
            14'b10_111111100101: DATA = 12'b100001010100;
            14'b10_111111100110: DATA = 12'b100001010001;
            14'b10_111111100111: DATA = 12'b100001001110;
            14'b10_111111101000: DATA = 12'b100001001011;
            14'b10_111111101001: DATA = 12'b100001001000;
            14'b10_111111101010: DATA = 12'b100001000101;
            14'b10_111111101011: DATA = 12'b100001000001;
            14'b10_111111101100: DATA = 12'b100000111110;
            14'b10_111111101101: DATA = 12'b100000111011;
            14'b10_111111101110: DATA = 12'b100000111000;
            14'b10_111111101111: DATA = 12'b100000110101;
            14'b10_111111110000: DATA = 12'b100000110010;
            14'b10_111111110001: DATA = 12'b100000101111;
            14'b10_111111110010: DATA = 12'b100000101011;
            14'b10_111111110011: DATA = 12'b100000101000;
            14'b10_111111110100: DATA = 12'b100000100101;
            14'b10_111111110101: DATA = 12'b100000100010;
            14'b10_111111110110: DATA = 12'b100000011111;
            14'b10_111111110111: DATA = 12'b100000011100;
            14'b10_111111111000: DATA = 12'b100000011001;
            14'b10_111111111001: DATA = 12'b100000010101;
            14'b10_111111111010: DATA = 12'b100000010010;
            14'b10_111111111011: DATA = 12'b100000001111;
            14'b10_111111111100: DATA = 12'b100000001100;
            14'b10_111111111101: DATA = 12'b100000001001;
            14'b10_111111111110: DATA = 12'b100000000110;
            14'b10_111111111111: DATA = 12'b100000000011;
            14'b11_000000000000: DATA = 12'b100000000000;
            14'b11_000000000001: DATA = 12'b100000000011;
            14'b11_000000000010: DATA = 12'b100000000110;
            14'b11_000000000011: DATA = 12'b100000001001;
            14'b11_000000000100: DATA = 12'b100000001100;
            14'b11_000000000101: DATA = 12'b100000001111;
            14'b11_000000000110: DATA = 12'b100000010010;
            14'b11_000000000111: DATA = 12'b100000010101;
            14'b11_000000001000: DATA = 12'b100000011001;
            14'b11_000000001001: DATA = 12'b100000011100;
            14'b11_000000001010: DATA = 12'b100000011111;
            14'b11_000000001011: DATA = 12'b100000100010;
            14'b11_000000001100: DATA = 12'b100000100101;
            14'b11_000000001101: DATA = 12'b100000101000;
            14'b11_000000001110: DATA = 12'b100000101011;
            14'b11_000000001111: DATA = 12'b100000101111;
            14'b11_000000010000: DATA = 12'b100000110010;
            14'b11_000000010001: DATA = 12'b100000110101;
            14'b11_000000010010: DATA = 12'b100000111000;
            14'b11_000000010011: DATA = 12'b100000111011;
            14'b11_000000010100: DATA = 12'b100000111110;
            14'b11_000000010101: DATA = 12'b100001000001;
            14'b11_000000010110: DATA = 12'b100001000101;
            14'b11_000000010111: DATA = 12'b100001001000;
            14'b11_000000011000: DATA = 12'b100001001011;
            14'b11_000000011001: DATA = 12'b100001001110;
            14'b11_000000011010: DATA = 12'b100001010001;
            14'b11_000000011011: DATA = 12'b100001010100;
            14'b11_000000011100: DATA = 12'b100001010111;
            14'b11_000000011101: DATA = 12'b100001011011;
            14'b11_000000011110: DATA = 12'b100001011110;
            14'b11_000000011111: DATA = 12'b100001100001;
            14'b11_000000100000: DATA = 12'b100001100100;
            14'b11_000000100001: DATA = 12'b100001100111;
            14'b11_000000100010: DATA = 12'b100001101010;
            14'b11_000000100011: DATA = 12'b100001101101;
            14'b11_000000100100: DATA = 12'b100001110000;
            14'b11_000000100101: DATA = 12'b100001110100;
            14'b11_000000100110: DATA = 12'b100001110111;
            14'b11_000000100111: DATA = 12'b100001111010;
            14'b11_000000101000: DATA = 12'b100001111101;
            14'b11_000000101001: DATA = 12'b100010000000;
            14'b11_000000101010: DATA = 12'b100010000011;
            14'b11_000000101011: DATA = 12'b100010000110;
            14'b11_000000101100: DATA = 12'b100010001010;
            14'b11_000000101101: DATA = 12'b100010001101;
            14'b11_000000101110: DATA = 12'b100010010000;
            14'b11_000000101111: DATA = 12'b100010010011;
            14'b11_000000110000: DATA = 12'b100010010110;
            14'b11_000000110001: DATA = 12'b100010011001;
            14'b11_000000110010: DATA = 12'b100010011100;
            14'b11_000000110011: DATA = 12'b100010011111;
            14'b11_000000110100: DATA = 12'b100010100011;
            14'b11_000000110101: DATA = 12'b100010100110;
            14'b11_000000110110: DATA = 12'b100010101001;
            14'b11_000000110111: DATA = 12'b100010101100;
            14'b11_000000111000: DATA = 12'b100010101111;
            14'b11_000000111001: DATA = 12'b100010110010;
            14'b11_000000111010: DATA = 12'b100010110101;
            14'b11_000000111011: DATA = 12'b100010111001;
            14'b11_000000111100: DATA = 12'b100010111100;
            14'b11_000000111101: DATA = 12'b100010111111;
            14'b11_000000111110: DATA = 12'b100011000010;
            14'b11_000000111111: DATA = 12'b100011000101;
            14'b11_000001000000: DATA = 12'b100011001000;
            14'b11_000001000001: DATA = 12'b100011001011;
            14'b11_000001000010: DATA = 12'b100011001110;
            14'b11_000001000011: DATA = 12'b100011010010;
            14'b11_000001000100: DATA = 12'b100011010101;
            14'b11_000001000101: DATA = 12'b100011011000;
            14'b11_000001000110: DATA = 12'b100011011011;
            14'b11_000001000111: DATA = 12'b100011011110;
            14'b11_000001001000: DATA = 12'b100011100001;
            14'b11_000001001001: DATA = 12'b100011100100;
            14'b11_000001001010: DATA = 12'b100011100111;
            14'b11_000001001011: DATA = 12'b100011101010;
            14'b11_000001001100: DATA = 12'b100011101110;
            14'b11_000001001101: DATA = 12'b100011110001;
            14'b11_000001001110: DATA = 12'b100011110100;
            14'b11_000001001111: DATA = 12'b100011110111;
            14'b11_000001010000: DATA = 12'b100011111010;
            14'b11_000001010001: DATA = 12'b100011111101;
            14'b11_000001010010: DATA = 12'b100100000000;
            14'b11_000001010011: DATA = 12'b100100000011;
            14'b11_000001010100: DATA = 12'b100100000111;
            14'b11_000001010101: DATA = 12'b100100001010;
            14'b11_000001010110: DATA = 12'b100100001101;
            14'b11_000001010111: DATA = 12'b100100010000;
            14'b11_000001011000: DATA = 12'b100100010011;
            14'b11_000001011001: DATA = 12'b100100010110;
            14'b11_000001011010: DATA = 12'b100100011001;
            14'b11_000001011011: DATA = 12'b100100011100;
            14'b11_000001011100: DATA = 12'b100100011111;
            14'b11_000001011101: DATA = 12'b100100100011;
            14'b11_000001011110: DATA = 12'b100100100110;
            14'b11_000001011111: DATA = 12'b100100101001;
            14'b11_000001100000: DATA = 12'b100100101100;
            14'b11_000001100001: DATA = 12'b100100101111;
            14'b11_000001100010: DATA = 12'b100100110010;
            14'b11_000001100011: DATA = 12'b100100110101;
            14'b11_000001100100: DATA = 12'b100100111000;
            14'b11_000001100101: DATA = 12'b100100111011;
            14'b11_000001100110: DATA = 12'b100100111110;
            14'b11_000001100111: DATA = 12'b100101000010;
            14'b11_000001101000: DATA = 12'b100101000101;
            14'b11_000001101001: DATA = 12'b100101001000;
            14'b11_000001101010: DATA = 12'b100101001011;
            14'b11_000001101011: DATA = 12'b100101001110;
            14'b11_000001101100: DATA = 12'b100101010001;
            14'b11_000001101101: DATA = 12'b100101010100;
            14'b11_000001101110: DATA = 12'b100101010111;
            14'b11_000001101111: DATA = 12'b100101011010;
            14'b11_000001110000: DATA = 12'b100101011101;
            14'b11_000001110001: DATA = 12'b100101100001;
            14'b11_000001110010: DATA = 12'b100101100100;
            14'b11_000001110011: DATA = 12'b100101100111;
            14'b11_000001110100: DATA = 12'b100101101010;
            14'b11_000001110101: DATA = 12'b100101101101;
            14'b11_000001110110: DATA = 12'b100101110000;
            14'b11_000001110111: DATA = 12'b100101110011;
            14'b11_000001111000: DATA = 12'b100101110110;
            14'b11_000001111001: DATA = 12'b100101111001;
            14'b11_000001111010: DATA = 12'b100101111100;
            14'b11_000001111011: DATA = 12'b100101111111;
            14'b11_000001111100: DATA = 12'b100110000011;
            14'b11_000001111101: DATA = 12'b100110000110;
            14'b11_000001111110: DATA = 12'b100110001001;
            14'b11_000001111111: DATA = 12'b100110001100;
            14'b11_000010000000: DATA = 12'b100110001111;
            14'b11_000010000001: DATA = 12'b100110010010;
            14'b11_000010000010: DATA = 12'b100110010101;
            14'b11_000010000011: DATA = 12'b100110011000;
            14'b11_000010000100: DATA = 12'b100110011011;
            14'b11_000010000101: DATA = 12'b100110011110;
            14'b11_000010000110: DATA = 12'b100110100001;
            14'b11_000010000111: DATA = 12'b100110100100;
            14'b11_000010001000: DATA = 12'b100110100111;
            14'b11_000010001001: DATA = 12'b100110101011;
            14'b11_000010001010: DATA = 12'b100110101110;
            14'b11_000010001011: DATA = 12'b100110110001;
            14'b11_000010001100: DATA = 12'b100110110100;
            14'b11_000010001101: DATA = 12'b100110110111;
            14'b11_000010001110: DATA = 12'b100110111010;
            14'b11_000010001111: DATA = 12'b100110111101;
            14'b11_000010010000: DATA = 12'b100111000000;
            14'b11_000010010001: DATA = 12'b100111000011;
            14'b11_000010010010: DATA = 12'b100111000110;
            14'b11_000010010011: DATA = 12'b100111001001;
            14'b11_000010010100: DATA = 12'b100111001100;
            14'b11_000010010101: DATA = 12'b100111001111;
            14'b11_000010010110: DATA = 12'b100111010010;
            14'b11_000010010111: DATA = 12'b100111010101;
            14'b11_000010011000: DATA = 12'b100111011000;
            14'b11_000010011001: DATA = 12'b100111011100;
            14'b11_000010011010: DATA = 12'b100111011111;
            14'b11_000010011011: DATA = 12'b100111100010;
            14'b11_000010011100: DATA = 12'b100111100101;
            14'b11_000010011101: DATA = 12'b100111101000;
            14'b11_000010011110: DATA = 12'b100111101011;
            14'b11_000010011111: DATA = 12'b100111101110;
            14'b11_000010100000: DATA = 12'b100111110001;
            14'b11_000010100001: DATA = 12'b100111110100;
            14'b11_000010100010: DATA = 12'b100111110111;
            14'b11_000010100011: DATA = 12'b100111111010;
            14'b11_000010100100: DATA = 12'b100111111101;
            14'b11_000010100101: DATA = 12'b101000000000;
            14'b11_000010100110: DATA = 12'b101000000011;
            14'b11_000010100111: DATA = 12'b101000000110;
            14'b11_000010101000: DATA = 12'b101000001001;
            14'b11_000010101001: DATA = 12'b101000001100;
            14'b11_000010101010: DATA = 12'b101000001111;
            14'b11_000010101011: DATA = 12'b101000010010;
            14'b11_000010101100: DATA = 12'b101000010101;
            14'b11_000010101101: DATA = 12'b101000011000;
            14'b11_000010101110: DATA = 12'b101000011011;
            14'b11_000010101111: DATA = 12'b101000011110;
            14'b11_000010110000: DATA = 12'b101000100001;
            14'b11_000010110001: DATA = 12'b101000100100;
            14'b11_000010110010: DATA = 12'b101000101000;
            14'b11_000010110011: DATA = 12'b101000101011;
            14'b11_000010110100: DATA = 12'b101000101110;
            14'b11_000010110101: DATA = 12'b101000110001;
            14'b11_000010110110: DATA = 12'b101000110100;
            14'b11_000010110111: DATA = 12'b101000110111;
            14'b11_000010111000: DATA = 12'b101000111010;
            14'b11_000010111001: DATA = 12'b101000111101;
            14'b11_000010111010: DATA = 12'b101001000000;
            14'b11_000010111011: DATA = 12'b101001000011;
            14'b11_000010111100: DATA = 12'b101001000110;
            14'b11_000010111101: DATA = 12'b101001001001;
            14'b11_000010111110: DATA = 12'b101001001100;
            14'b11_000010111111: DATA = 12'b101001001111;
            14'b11_000011000000: DATA = 12'b101001010010;
            14'b11_000011000001: DATA = 12'b101001010101;
            14'b11_000011000010: DATA = 12'b101001011000;
            14'b11_000011000011: DATA = 12'b101001011011;
            14'b11_000011000100: DATA = 12'b101001011110;
            14'b11_000011000101: DATA = 12'b101001100001;
            14'b11_000011000110: DATA = 12'b101001100100;
            14'b11_000011000111: DATA = 12'b101001100111;
            14'b11_000011001000: DATA = 12'b101001101010;
            14'b11_000011001001: DATA = 12'b101001101101;
            14'b11_000011001010: DATA = 12'b101001110000;
            14'b11_000011001011: DATA = 12'b101001110011;
            14'b11_000011001100: DATA = 12'b101001110110;
            14'b11_000011001101: DATA = 12'b101001111001;
            14'b11_000011001110: DATA = 12'b101001111100;
            14'b11_000011001111: DATA = 12'b101001111111;
            14'b11_000011010000: DATA = 12'b101010000010;
            14'b11_000011010001: DATA = 12'b101010000101;
            14'b11_000011010010: DATA = 12'b101010001000;
            14'b11_000011010011: DATA = 12'b101010001011;
            14'b11_000011010100: DATA = 12'b101010001110;
            14'b11_000011010101: DATA = 12'b101010010000;
            14'b11_000011010110: DATA = 12'b101010010011;
            14'b11_000011010111: DATA = 12'b101010010110;
            14'b11_000011011000: DATA = 12'b101010011001;
            14'b11_000011011001: DATA = 12'b101010011100;
            14'b11_000011011010: DATA = 12'b101010011111;
            14'b11_000011011011: DATA = 12'b101010100010;
            14'b11_000011011100: DATA = 12'b101010100101;
            14'b11_000011011101: DATA = 12'b101010101000;
            14'b11_000011011110: DATA = 12'b101010101011;
            14'b11_000011011111: DATA = 12'b101010101110;
            14'b11_000011100000: DATA = 12'b101010110001;
            14'b11_000011100001: DATA = 12'b101010110100;
            14'b11_000011100010: DATA = 12'b101010110111;
            14'b11_000011100011: DATA = 12'b101010111010;
            14'b11_000011100100: DATA = 12'b101010111101;
            14'b11_000011100101: DATA = 12'b101011000000;
            14'b11_000011100110: DATA = 12'b101011000011;
            14'b11_000011100111: DATA = 12'b101011000110;
            14'b11_000011101000: DATA = 12'b101011001001;
            14'b11_000011101001: DATA = 12'b101011001100;
            14'b11_000011101010: DATA = 12'b101011001111;
            14'b11_000011101011: DATA = 12'b101011010010;
            14'b11_000011101100: DATA = 12'b101011010100;
            14'b11_000011101101: DATA = 12'b101011010111;
            14'b11_000011101110: DATA = 12'b101011011010;
            14'b11_000011101111: DATA = 12'b101011011101;
            14'b11_000011110000: DATA = 12'b101011100000;
            14'b11_000011110001: DATA = 12'b101011100011;
            14'b11_000011110010: DATA = 12'b101011100110;
            14'b11_000011110011: DATA = 12'b101011101001;
            14'b11_000011110100: DATA = 12'b101011101100;
            14'b11_000011110101: DATA = 12'b101011101111;
            14'b11_000011110110: DATA = 12'b101011110010;
            14'b11_000011110111: DATA = 12'b101011110101;
            14'b11_000011111000: DATA = 12'b101011111000;
            14'b11_000011111001: DATA = 12'b101011111011;
            14'b11_000011111010: DATA = 12'b101011111101;
            14'b11_000011111011: DATA = 12'b101100000000;
            14'b11_000011111100: DATA = 12'b101100000011;
            14'b11_000011111101: DATA = 12'b101100000110;
            14'b11_000011111110: DATA = 12'b101100001001;
            14'b11_000011111111: DATA = 12'b101100001100;
            14'b11_000100000000: DATA = 12'b101100001111;
            14'b11_000100000001: DATA = 12'b101100010010;
            14'b11_000100000010: DATA = 12'b101100010101;
            14'b11_000100000011: DATA = 12'b101100011000;
            14'b11_000100000100: DATA = 12'b101100011010;
            14'b11_000100000101: DATA = 12'b101100011101;
            14'b11_000100000110: DATA = 12'b101100100000;
            14'b11_000100000111: DATA = 12'b101100100011;
            14'b11_000100001000: DATA = 12'b101100100110;
            14'b11_000100001001: DATA = 12'b101100101001;
            14'b11_000100001010: DATA = 12'b101100101100;
            14'b11_000100001011: DATA = 12'b101100101111;
            14'b11_000100001100: DATA = 12'b101100110010;
            14'b11_000100001101: DATA = 12'b101100110100;
            14'b11_000100001110: DATA = 12'b101100110111;
            14'b11_000100001111: DATA = 12'b101100111010;
            14'b11_000100010000: DATA = 12'b101100111101;
            14'b11_000100010001: DATA = 12'b101101000000;
            14'b11_000100010010: DATA = 12'b101101000011;
            14'b11_000100010011: DATA = 12'b101101000110;
            14'b11_000100010100: DATA = 12'b101101001000;
            14'b11_000100010101: DATA = 12'b101101001011;
            14'b11_000100010110: DATA = 12'b101101001110;
            14'b11_000100010111: DATA = 12'b101101010001;
            14'b11_000100011000: DATA = 12'b101101010100;
            14'b11_000100011001: DATA = 12'b101101010111;
            14'b11_000100011010: DATA = 12'b101101011010;
            14'b11_000100011011: DATA = 12'b101101011100;
            14'b11_000100011100: DATA = 12'b101101011111;
            14'b11_000100011101: DATA = 12'b101101100010;
            14'b11_000100011110: DATA = 12'b101101100101;
            14'b11_000100011111: DATA = 12'b101101101000;
            14'b11_000100100000: DATA = 12'b101101101011;
            14'b11_000100100001: DATA = 12'b101101101110;
            14'b11_000100100010: DATA = 12'b101101110000;
            14'b11_000100100011: DATA = 12'b101101110011;
            14'b11_000100100100: DATA = 12'b101101110110;
            14'b11_000100100101: DATA = 12'b101101111001;
            14'b11_000100100110: DATA = 12'b101101111100;
            14'b11_000100100111: DATA = 12'b101101111111;
            14'b11_000100101000: DATA = 12'b101110000001;
            14'b11_000100101001: DATA = 12'b101110000100;
            14'b11_000100101010: DATA = 12'b101110000111;
            14'b11_000100101011: DATA = 12'b101110001010;
            14'b11_000100101100: DATA = 12'b101110001101;
            14'b11_000100101101: DATA = 12'b101110001111;
            14'b11_000100101110: DATA = 12'b101110010010;
            14'b11_000100101111: DATA = 12'b101110010101;
            14'b11_000100110000: DATA = 12'b101110011000;
            14'b11_000100110001: DATA = 12'b101110011011;
            14'b11_000100110010: DATA = 12'b101110011101;
            14'b11_000100110011: DATA = 12'b101110100000;
            14'b11_000100110100: DATA = 12'b101110100011;
            14'b11_000100110101: DATA = 12'b101110100110;
            14'b11_000100110110: DATA = 12'b101110101001;
            14'b11_000100110111: DATA = 12'b101110101011;
            14'b11_000100111000: DATA = 12'b101110101110;
            14'b11_000100111001: DATA = 12'b101110110001;
            14'b11_000100111010: DATA = 12'b101110110100;
            14'b11_000100111011: DATA = 12'b101110110111;
            14'b11_000100111100: DATA = 12'b101110111001;
            14'b11_000100111101: DATA = 12'b101110111100;
            14'b11_000100111110: DATA = 12'b101110111111;
            14'b11_000100111111: DATA = 12'b101111000010;
            14'b11_000101000000: DATA = 12'b101111000100;
            14'b11_000101000001: DATA = 12'b101111000111;
            14'b11_000101000010: DATA = 12'b101111001010;
            14'b11_000101000011: DATA = 12'b101111001101;
            14'b11_000101000100: DATA = 12'b101111010000;
            14'b11_000101000101: DATA = 12'b101111010010;
            14'b11_000101000110: DATA = 12'b101111010101;
            14'b11_000101000111: DATA = 12'b101111011000;
            14'b11_000101001000: DATA = 12'b101111011011;
            14'b11_000101001001: DATA = 12'b101111011101;
            14'b11_000101001010: DATA = 12'b101111100000;
            14'b11_000101001011: DATA = 12'b101111100011;
            14'b11_000101001100: DATA = 12'b101111100110;
            14'b11_000101001101: DATA = 12'b101111101000;
            14'b11_000101001110: DATA = 12'b101111101011;
            14'b11_000101001111: DATA = 12'b101111101110;
            14'b11_000101010000: DATA = 12'b101111110000;
            14'b11_000101010001: DATA = 12'b101111110011;
            14'b11_000101010010: DATA = 12'b101111110110;
            14'b11_000101010011: DATA = 12'b101111111001;
            14'b11_000101010100: DATA = 12'b101111111011;
            14'b11_000101010101: DATA = 12'b101111111110;
            14'b11_000101010110: DATA = 12'b110000000001;
            14'b11_000101010111: DATA = 12'b110000000100;
            14'b11_000101011000: DATA = 12'b110000000110;
            14'b11_000101011001: DATA = 12'b110000001001;
            14'b11_000101011010: DATA = 12'b110000001100;
            14'b11_000101011011: DATA = 12'b110000001110;
            14'b11_000101011100: DATA = 12'b110000010001;
            14'b11_000101011101: DATA = 12'b110000010100;
            14'b11_000101011110: DATA = 12'b110000010110;
            14'b11_000101011111: DATA = 12'b110000011001;
            14'b11_000101100000: DATA = 12'b110000011100;
            14'b11_000101100001: DATA = 12'b110000011111;
            14'b11_000101100010: DATA = 12'b110000100001;
            14'b11_000101100011: DATA = 12'b110000100100;
            14'b11_000101100100: DATA = 12'b110000100111;
            14'b11_000101100101: DATA = 12'b110000101001;
            14'b11_000101100110: DATA = 12'b110000101100;
            14'b11_000101100111: DATA = 12'b110000101111;
            14'b11_000101101000: DATA = 12'b110000110001;
            14'b11_000101101001: DATA = 12'b110000110100;
            14'b11_000101101010: DATA = 12'b110000110111;
            14'b11_000101101011: DATA = 12'b110000111001;
            14'b11_000101101100: DATA = 12'b110000111100;
            14'b11_000101101101: DATA = 12'b110000111111;
            14'b11_000101101110: DATA = 12'b110001000001;
            14'b11_000101101111: DATA = 12'b110001000100;
            14'b11_000101110000: DATA = 12'b110001000111;
            14'b11_000101110001: DATA = 12'b110001001001;
            14'b11_000101110010: DATA = 12'b110001001100;
            14'b11_000101110011: DATA = 12'b110001001111;
            14'b11_000101110100: DATA = 12'b110001010001;
            14'b11_000101110101: DATA = 12'b110001010100;
            14'b11_000101110110: DATA = 12'b110001010111;
            14'b11_000101110111: DATA = 12'b110001011001;
            14'b11_000101111000: DATA = 12'b110001011100;
            14'b11_000101111001: DATA = 12'b110001011110;
            14'b11_000101111010: DATA = 12'b110001100001;
            14'b11_000101111011: DATA = 12'b110001100100;
            14'b11_000101111100: DATA = 12'b110001100110;
            14'b11_000101111101: DATA = 12'b110001101001;
            14'b11_000101111110: DATA = 12'b110001101100;
            14'b11_000101111111: DATA = 12'b110001101110;
            14'b11_000110000000: DATA = 12'b110001110001;
            14'b11_000110000001: DATA = 12'b110001110011;
            14'b11_000110000010: DATA = 12'b110001110110;
            14'b11_000110000011: DATA = 12'b110001111001;
            14'b11_000110000100: DATA = 12'b110001111011;
            14'b11_000110000101: DATA = 12'b110001111110;
            14'b11_000110000110: DATA = 12'b110010000000;
            14'b11_000110000111: DATA = 12'b110010000011;
            14'b11_000110001000: DATA = 12'b110010000110;
            14'b11_000110001001: DATA = 12'b110010001000;
            14'b11_000110001010: DATA = 12'b110010001011;
            14'b11_000110001011: DATA = 12'b110010001101;
            14'b11_000110001100: DATA = 12'b110010010000;
            14'b11_000110001101: DATA = 12'b110010010010;
            14'b11_000110001110: DATA = 12'b110010010101;
            14'b11_000110001111: DATA = 12'b110010011000;
            14'b11_000110010000: DATA = 12'b110010011010;
            14'b11_000110010001: DATA = 12'b110010011101;
            14'b11_000110010010: DATA = 12'b110010011111;
            14'b11_000110010011: DATA = 12'b110010100010;
            14'b11_000110010100: DATA = 12'b110010100100;
            14'b11_000110010101: DATA = 12'b110010100111;
            14'b11_000110010110: DATA = 12'b110010101010;
            14'b11_000110010111: DATA = 12'b110010101100;
            14'b11_000110011000: DATA = 12'b110010101111;
            14'b11_000110011001: DATA = 12'b110010110001;
            14'b11_000110011010: DATA = 12'b110010110100;
            14'b11_000110011011: DATA = 12'b110010110110;
            14'b11_000110011100: DATA = 12'b110010111001;
            14'b11_000110011101: DATA = 12'b110010111011;
            14'b11_000110011110: DATA = 12'b110010111110;
            14'b11_000110011111: DATA = 12'b110011000000;
            14'b11_000110100000: DATA = 12'b110011000011;
            14'b11_000110100001: DATA = 12'b110011000101;
            14'b11_000110100010: DATA = 12'b110011001000;
            14'b11_000110100011: DATA = 12'b110011001010;
            14'b11_000110100100: DATA = 12'b110011001101;
            14'b11_000110100101: DATA = 12'b110011001111;
            14'b11_000110100110: DATA = 12'b110011010010;
            14'b11_000110100111: DATA = 12'b110011010100;
            14'b11_000110101000: DATA = 12'b110011010111;
            14'b11_000110101001: DATA = 12'b110011011001;
            14'b11_000110101010: DATA = 12'b110011011100;
            14'b11_000110101011: DATA = 12'b110011011110;
            14'b11_000110101100: DATA = 12'b110011100001;
            14'b11_000110101101: DATA = 12'b110011100011;
            14'b11_000110101110: DATA = 12'b110011100110;
            14'b11_000110101111: DATA = 12'b110011101000;
            14'b11_000110110000: DATA = 12'b110011101011;
            14'b11_000110110001: DATA = 12'b110011101101;
            14'b11_000110110010: DATA = 12'b110011110000;
            14'b11_000110110011: DATA = 12'b110011110010;
            14'b11_000110110100: DATA = 12'b110011110101;
            14'b11_000110110101: DATA = 12'b110011110111;
            14'b11_000110110110: DATA = 12'b110011111010;
            14'b11_000110110111: DATA = 12'b110011111100;
            14'b11_000110111000: DATA = 12'b110011111111;
            14'b11_000110111001: DATA = 12'b110100000001;
            14'b11_000110111010: DATA = 12'b110100000011;
            14'b11_000110111011: DATA = 12'b110100000110;
            14'b11_000110111100: DATA = 12'b110100001000;
            14'b11_000110111101: DATA = 12'b110100001011;
            14'b11_000110111110: DATA = 12'b110100001101;
            14'b11_000110111111: DATA = 12'b110100010000;
            14'b11_000111000000: DATA = 12'b110100010010;
            14'b11_000111000001: DATA = 12'b110100010101;
            14'b11_000111000010: DATA = 12'b110100010111;
            14'b11_000111000011: DATA = 12'b110100011001;
            14'b11_000111000100: DATA = 12'b110100011100;
            14'b11_000111000101: DATA = 12'b110100011110;
            14'b11_000111000110: DATA = 12'b110100100001;
            14'b11_000111000111: DATA = 12'b110100100011;
            14'b11_000111001000: DATA = 12'b110100100101;
            14'b11_000111001001: DATA = 12'b110100101000;
            14'b11_000111001010: DATA = 12'b110100101010;
            14'b11_000111001011: DATA = 12'b110100101101;
            14'b11_000111001100: DATA = 12'b110100101111;
            14'b11_000111001101: DATA = 12'b110100110001;
            14'b11_000111001110: DATA = 12'b110100110100;
            14'b11_000111001111: DATA = 12'b110100110110;
            14'b11_000111010000: DATA = 12'b110100111001;
            14'b11_000111010001: DATA = 12'b110100111011;
            14'b11_000111010010: DATA = 12'b110100111101;
            14'b11_000111010011: DATA = 12'b110101000000;
            14'b11_000111010100: DATA = 12'b110101000010;
            14'b11_000111010101: DATA = 12'b110101000100;
            14'b11_000111010110: DATA = 12'b110101000111;
            14'b11_000111010111: DATA = 12'b110101001001;
            14'b11_000111011000: DATA = 12'b110101001011;
            14'b11_000111011001: DATA = 12'b110101001110;
            14'b11_000111011010: DATA = 12'b110101010000;
            14'b11_000111011011: DATA = 12'b110101010011;
            14'b11_000111011100: DATA = 12'b110101010101;
            14'b11_000111011101: DATA = 12'b110101010111;
            14'b11_000111011110: DATA = 12'b110101011010;
            14'b11_000111011111: DATA = 12'b110101011100;
            14'b11_000111100000: DATA = 12'b110101011110;
            14'b11_000111100001: DATA = 12'b110101100001;
            14'b11_000111100010: DATA = 12'b110101100011;
            14'b11_000111100011: DATA = 12'b110101100101;
            14'b11_000111100100: DATA = 12'b110101100111;
            14'b11_000111100101: DATA = 12'b110101101010;
            14'b11_000111100110: DATA = 12'b110101101100;
            14'b11_000111100111: DATA = 12'b110101101110;
            14'b11_000111101000: DATA = 12'b110101110001;
            14'b11_000111101001: DATA = 12'b110101110011;
            14'b11_000111101010: DATA = 12'b110101110101;
            14'b11_000111101011: DATA = 12'b110101111000;
            14'b11_000111101100: DATA = 12'b110101111010;
            14'b11_000111101101: DATA = 12'b110101111100;
            14'b11_000111101110: DATA = 12'b110101111110;
            14'b11_000111101111: DATA = 12'b110110000001;
            14'b11_000111110000: DATA = 12'b110110000011;
            14'b11_000111110001: DATA = 12'b110110000101;
            14'b11_000111110010: DATA = 12'b110110001000;
            14'b11_000111110011: DATA = 12'b110110001010;
            14'b11_000111110100: DATA = 12'b110110001100;
            14'b11_000111110101: DATA = 12'b110110001110;
            14'b11_000111110110: DATA = 12'b110110010001;
            14'b11_000111110111: DATA = 12'b110110010011;
            14'b11_000111111000: DATA = 12'b110110010101;
            14'b11_000111111001: DATA = 12'b110110010111;
            14'b11_000111111010: DATA = 12'b110110011010;
            14'b11_000111111011: DATA = 12'b110110011100;
            14'b11_000111111100: DATA = 12'b110110011110;
            14'b11_000111111101: DATA = 12'b110110100000;
            14'b11_000111111110: DATA = 12'b110110100011;
            14'b11_000111111111: DATA = 12'b110110100101;
            14'b11_001000000000: DATA = 12'b110110100111;
            14'b11_001000000001: DATA = 12'b110110101001;
            14'b11_001000000010: DATA = 12'b110110101011;
            14'b11_001000000011: DATA = 12'b110110101110;
            14'b11_001000000100: DATA = 12'b110110110000;
            14'b11_001000000101: DATA = 12'b110110110010;
            14'b11_001000000110: DATA = 12'b110110110100;
            14'b11_001000000111: DATA = 12'b110110110110;
            14'b11_001000001000: DATA = 12'b110110111001;
            14'b11_001000001001: DATA = 12'b110110111011;
            14'b11_001000001010: DATA = 12'b110110111101;
            14'b11_001000001011: DATA = 12'b110110111111;
            14'b11_001000001100: DATA = 12'b110111000001;
            14'b11_001000001101: DATA = 12'b110111000100;
            14'b11_001000001110: DATA = 12'b110111000110;
            14'b11_001000001111: DATA = 12'b110111001000;
            14'b11_001000010000: DATA = 12'b110111001010;
            14'b11_001000010001: DATA = 12'b110111001100;
            14'b11_001000010010: DATA = 12'b110111001110;
            14'b11_001000010011: DATA = 12'b110111010001;
            14'b11_001000010100: DATA = 12'b110111010011;
            14'b11_001000010101: DATA = 12'b110111010101;
            14'b11_001000010110: DATA = 12'b110111010111;
            14'b11_001000010111: DATA = 12'b110111011001;
            14'b11_001000011000: DATA = 12'b110111011011;
            14'b11_001000011001: DATA = 12'b110111011101;
            14'b11_001000011010: DATA = 12'b110111100000;
            14'b11_001000011011: DATA = 12'b110111100010;
            14'b11_001000011100: DATA = 12'b110111100100;
            14'b11_001000011101: DATA = 12'b110111100110;
            14'b11_001000011110: DATA = 12'b110111101000;
            14'b11_001000011111: DATA = 12'b110111101010;
            14'b11_001000100000: DATA = 12'b110111101100;
            14'b11_001000100001: DATA = 12'b110111101110;
            14'b11_001000100010: DATA = 12'b110111110000;
            14'b11_001000100011: DATA = 12'b110111110011;
            14'b11_001000100100: DATA = 12'b110111110101;
            14'b11_001000100101: DATA = 12'b110111110111;
            14'b11_001000100110: DATA = 12'b110111111001;
            14'b11_001000100111: DATA = 12'b110111111011;
            14'b11_001000101000: DATA = 12'b110111111101;
            14'b11_001000101001: DATA = 12'b110111111111;
            14'b11_001000101010: DATA = 12'b111000000001;
            14'b11_001000101011: DATA = 12'b111000000011;
            14'b11_001000101100: DATA = 12'b111000000101;
            14'b11_001000101101: DATA = 12'b111000000111;
            14'b11_001000101110: DATA = 12'b111000001001;
            14'b11_001000101111: DATA = 12'b111000001011;
            14'b11_001000110000: DATA = 12'b111000001110;
            14'b11_001000110001: DATA = 12'b111000010000;
            14'b11_001000110010: DATA = 12'b111000010010;
            14'b11_001000110011: DATA = 12'b111000010100;
            14'b11_001000110100: DATA = 12'b111000010110;
            14'b11_001000110101: DATA = 12'b111000011000;
            14'b11_001000110110: DATA = 12'b111000011010;
            14'b11_001000110111: DATA = 12'b111000011100;
            14'b11_001000111000: DATA = 12'b111000011110;
            14'b11_001000111001: DATA = 12'b111000100000;
            14'b11_001000111010: DATA = 12'b111000100010;
            14'b11_001000111011: DATA = 12'b111000100100;
            14'b11_001000111100: DATA = 12'b111000100110;
            14'b11_001000111101: DATA = 12'b111000101000;
            14'b11_001000111110: DATA = 12'b111000101010;
            14'b11_001000111111: DATA = 12'b111000101100;
            14'b11_001001000000: DATA = 12'b111000101110;
            14'b11_001001000001: DATA = 12'b111000110000;
            14'b11_001001000010: DATA = 12'b111000110010;
            14'b11_001001000011: DATA = 12'b111000110100;
            14'b11_001001000100: DATA = 12'b111000110110;
            14'b11_001001000101: DATA = 12'b111000111000;
            14'b11_001001000110: DATA = 12'b111000111010;
            14'b11_001001000111: DATA = 12'b111000111100;
            14'b11_001001001000: DATA = 12'b111000111110;
            14'b11_001001001001: DATA = 12'b111001000000;
            14'b11_001001001010: DATA = 12'b111001000010;
            14'b11_001001001011: DATA = 12'b111001000100;
            14'b11_001001001100: DATA = 12'b111001000101;
            14'b11_001001001101: DATA = 12'b111001000111;
            14'b11_001001001110: DATA = 12'b111001001001;
            14'b11_001001001111: DATA = 12'b111001001011;
            14'b11_001001010000: DATA = 12'b111001001101;
            14'b11_001001010001: DATA = 12'b111001001111;
            14'b11_001001010010: DATA = 12'b111001010001;
            14'b11_001001010011: DATA = 12'b111001010011;
            14'b11_001001010100: DATA = 12'b111001010101;
            14'b11_001001010101: DATA = 12'b111001010111;
            14'b11_001001010110: DATA = 12'b111001011001;
            14'b11_001001010111: DATA = 12'b111001011011;
            14'b11_001001011000: DATA = 12'b111001011101;
            14'b11_001001011001: DATA = 12'b111001011110;
            14'b11_001001011010: DATA = 12'b111001100000;
            14'b11_001001011011: DATA = 12'b111001100010;
            14'b11_001001011100: DATA = 12'b111001100100;
            14'b11_001001011101: DATA = 12'b111001100110;
            14'b11_001001011110: DATA = 12'b111001101000;
            14'b11_001001011111: DATA = 12'b111001101010;
            14'b11_001001100000: DATA = 12'b111001101100;
            14'b11_001001100001: DATA = 12'b111001101110;
            14'b11_001001100010: DATA = 12'b111001101111;
            14'b11_001001100011: DATA = 12'b111001110001;
            14'b11_001001100100: DATA = 12'b111001110011;
            14'b11_001001100101: DATA = 12'b111001110101;
            14'b11_001001100110: DATA = 12'b111001110111;
            14'b11_001001100111: DATA = 12'b111001111001;
            14'b11_001001101000: DATA = 12'b111001111011;
            14'b11_001001101001: DATA = 12'b111001111100;
            14'b11_001001101010: DATA = 12'b111001111110;
            14'b11_001001101011: DATA = 12'b111010000000;
            14'b11_001001101100: DATA = 12'b111010000010;
            14'b11_001001101101: DATA = 12'b111010000100;
            14'b11_001001101110: DATA = 12'b111010000101;
            14'b11_001001101111: DATA = 12'b111010000111;
            14'b11_001001110000: DATA = 12'b111010001001;
            14'b11_001001110001: DATA = 12'b111010001011;
            14'b11_001001110010: DATA = 12'b111010001101;
            14'b11_001001110011: DATA = 12'b111010001111;
            14'b11_001001110100: DATA = 12'b111010010000;
            14'b11_001001110101: DATA = 12'b111010010010;
            14'b11_001001110110: DATA = 12'b111010010100;
            14'b11_001001110111: DATA = 12'b111010010110;
            14'b11_001001111000: DATA = 12'b111010010111;
            14'b11_001001111001: DATA = 12'b111010011001;
            14'b11_001001111010: DATA = 12'b111010011011;
            14'b11_001001111011: DATA = 12'b111010011101;
            14'b11_001001111100: DATA = 12'b111010011111;
            14'b11_001001111101: DATA = 12'b111010100000;
            14'b11_001001111110: DATA = 12'b111010100010;
            14'b11_001001111111: DATA = 12'b111010100100;
            14'b11_001010000000: DATA = 12'b111010100110;
            14'b11_001010000001: DATA = 12'b111010100111;
            14'b11_001010000010: DATA = 12'b111010101001;
            14'b11_001010000011: DATA = 12'b111010101011;
            14'b11_001010000100: DATA = 12'b111010101100;
            14'b11_001010000101: DATA = 12'b111010101110;
            14'b11_001010000110: DATA = 12'b111010110000;
            14'b11_001010000111: DATA = 12'b111010110010;
            14'b11_001010001000: DATA = 12'b111010110011;
            14'b11_001010001001: DATA = 12'b111010110101;
            14'b11_001010001010: DATA = 12'b111010110111;
            14'b11_001010001011: DATA = 12'b111010111000;
            14'b11_001010001100: DATA = 12'b111010111010;
            14'b11_001010001101: DATA = 12'b111010111100;
            14'b11_001010001110: DATA = 12'b111010111110;
            14'b11_001010001111: DATA = 12'b111010111111;
            14'b11_001010010000: DATA = 12'b111011000001;
            14'b11_001010010001: DATA = 12'b111011000011;
            14'b11_001010010010: DATA = 12'b111011000100;
            14'b11_001010010011: DATA = 12'b111011000110;
            14'b11_001010010100: DATA = 12'b111011001000;
            14'b11_001010010101: DATA = 12'b111011001001;
            14'b11_001010010110: DATA = 12'b111011001011;
            14'b11_001010010111: DATA = 12'b111011001101;
            14'b11_001010011000: DATA = 12'b111011001110;
            14'b11_001010011001: DATA = 12'b111011010000;
            14'b11_001010011010: DATA = 12'b111011010010;
            14'b11_001010011011: DATA = 12'b111011010011;
            14'b11_001010011100: DATA = 12'b111011010101;
            14'b11_001010011101: DATA = 12'b111011010110;
            14'b11_001010011110: DATA = 12'b111011011000;
            14'b11_001010011111: DATA = 12'b111011011010;
            14'b11_001010100000: DATA = 12'b111011011011;
            14'b11_001010100001: DATA = 12'b111011011101;
            14'b11_001010100010: DATA = 12'b111011011110;
            14'b11_001010100011: DATA = 12'b111011100000;
            14'b11_001010100100: DATA = 12'b111011100010;
            14'b11_001010100101: DATA = 12'b111011100011;
            14'b11_001010100110: DATA = 12'b111011100101;
            14'b11_001010100111: DATA = 12'b111011100110;
            14'b11_001010101000: DATA = 12'b111011101000;
            14'b11_001010101001: DATA = 12'b111011101010;
            14'b11_001010101010: DATA = 12'b111011101011;
            14'b11_001010101011: DATA = 12'b111011101101;
            14'b11_001010101100: DATA = 12'b111011101110;
            14'b11_001010101101: DATA = 12'b111011110000;
            14'b11_001010101110: DATA = 12'b111011110001;
            14'b11_001010101111: DATA = 12'b111011110011;
            14'b11_001010110000: DATA = 12'b111011110101;
            14'b11_001010110001: DATA = 12'b111011110110;
            14'b11_001010110010: DATA = 12'b111011111000;
            14'b11_001010110011: DATA = 12'b111011111001;
            14'b11_001010110100: DATA = 12'b111011111011;
            14'b11_001010110101: DATA = 12'b111011111100;
            14'b11_001010110110: DATA = 12'b111011111110;
            14'b11_001010110111: DATA = 12'b111011111111;
            14'b11_001010111000: DATA = 12'b111100000001;
            14'b11_001010111001: DATA = 12'b111100000010;
            14'b11_001010111010: DATA = 12'b111100000100;
            14'b11_001010111011: DATA = 12'b111100000101;
            14'b11_001010111100: DATA = 12'b111100000111;
            14'b11_001010111101: DATA = 12'b111100001000;
            14'b11_001010111110: DATA = 12'b111100001010;
            14'b11_001010111111: DATA = 12'b111100001011;
            14'b11_001011000000: DATA = 12'b111100001101;
            14'b11_001011000001: DATA = 12'b111100001110;
            14'b11_001011000010: DATA = 12'b111100010000;
            14'b11_001011000011: DATA = 12'b111100010001;
            14'b11_001011000100: DATA = 12'b111100010011;
            14'b11_001011000101: DATA = 12'b111100010100;
            14'b11_001011000110: DATA = 12'b111100010110;
            14'b11_001011000111: DATA = 12'b111100010111;
            14'b11_001011001000: DATA = 12'b111100011000;
            14'b11_001011001001: DATA = 12'b111100011010;
            14'b11_001011001010: DATA = 12'b111100011011;
            14'b11_001011001011: DATA = 12'b111100011101;
            14'b11_001011001100: DATA = 12'b111100011110;
            14'b11_001011001101: DATA = 12'b111100100000;
            14'b11_001011001110: DATA = 12'b111100100001;
            14'b11_001011001111: DATA = 12'b111100100011;
            14'b11_001011010000: DATA = 12'b111100100100;
            14'b11_001011010001: DATA = 12'b111100100101;
            14'b11_001011010010: DATA = 12'b111100100111;
            14'b11_001011010011: DATA = 12'b111100101000;
            14'b11_001011010100: DATA = 12'b111100101010;
            14'b11_001011010101: DATA = 12'b111100101011;
            14'b11_001011010110: DATA = 12'b111100101100;
            14'b11_001011010111: DATA = 12'b111100101110;
            14'b11_001011011000: DATA = 12'b111100101111;
            14'b11_001011011001: DATA = 12'b111100110000;
            14'b11_001011011010: DATA = 12'b111100110010;
            14'b11_001011011011: DATA = 12'b111100110011;
            14'b11_001011011100: DATA = 12'b111100110101;
            14'b11_001011011101: DATA = 12'b111100110110;
            14'b11_001011011110: DATA = 12'b111100110111;
            14'b11_001011011111: DATA = 12'b111100111001;
            14'b11_001011100000: DATA = 12'b111100111010;
            14'b11_001011100001: DATA = 12'b111100111011;
            14'b11_001011100010: DATA = 12'b111100111101;
            14'b11_001011100011: DATA = 12'b111100111110;
            14'b11_001011100100: DATA = 12'b111100111111;
            14'b11_001011100101: DATA = 12'b111101000001;
            14'b11_001011100110: DATA = 12'b111101000010;
            14'b11_001011100111: DATA = 12'b111101000011;
            14'b11_001011101000: DATA = 12'b111101000101;
            14'b11_001011101001: DATA = 12'b111101000110;
            14'b11_001011101010: DATA = 12'b111101000111;
            14'b11_001011101011: DATA = 12'b111101001000;
            14'b11_001011101100: DATA = 12'b111101001010;
            14'b11_001011101101: DATA = 12'b111101001011;
            14'b11_001011101110: DATA = 12'b111101001100;
            14'b11_001011101111: DATA = 12'b111101001110;
            14'b11_001011110000: DATA = 12'b111101001111;
            14'b11_001011110001: DATA = 12'b111101010000;
            14'b11_001011110010: DATA = 12'b111101010001;
            14'b11_001011110011: DATA = 12'b111101010011;
            14'b11_001011110100: DATA = 12'b111101010100;
            14'b11_001011110101: DATA = 12'b111101010101;
            14'b11_001011110110: DATA = 12'b111101010110;
            14'b11_001011110111: DATA = 12'b111101011000;
            14'b11_001011111000: DATA = 12'b111101011001;
            14'b11_001011111001: DATA = 12'b111101011010;
            14'b11_001011111010: DATA = 12'b111101011011;
            14'b11_001011111011: DATA = 12'b111101011101;
            14'b11_001011111100: DATA = 12'b111101011110;
            14'b11_001011111101: DATA = 12'b111101011111;
            14'b11_001011111110: DATA = 12'b111101100000;
            14'b11_001011111111: DATA = 12'b111101100001;
            14'b11_001100000000: DATA = 12'b111101100011;
            14'b11_001100000001: DATA = 12'b111101100100;
            14'b11_001100000010: DATA = 12'b111101100101;
            14'b11_001100000011: DATA = 12'b111101100110;
            14'b11_001100000100: DATA = 12'b111101100111;
            14'b11_001100000101: DATA = 12'b111101101001;
            14'b11_001100000110: DATA = 12'b111101101010;
            14'b11_001100000111: DATA = 12'b111101101011;
            14'b11_001100001000: DATA = 12'b111101101100;
            14'b11_001100001001: DATA = 12'b111101101101;
            14'b11_001100001010: DATA = 12'b111101101110;
            14'b11_001100001011: DATA = 12'b111101110000;
            14'b11_001100001100: DATA = 12'b111101110001;
            14'b11_001100001101: DATA = 12'b111101110010;
            14'b11_001100001110: DATA = 12'b111101110011;
            14'b11_001100001111: DATA = 12'b111101110100;
            14'b11_001100010000: DATA = 12'b111101110101;
            14'b11_001100010001: DATA = 12'b111101110110;
            14'b11_001100010010: DATA = 12'b111101111000;
            14'b11_001100010011: DATA = 12'b111101111001;
            14'b11_001100010100: DATA = 12'b111101111010;
            14'b11_001100010101: DATA = 12'b111101111011;
            14'b11_001100010110: DATA = 12'b111101111100;
            14'b11_001100010111: DATA = 12'b111101111101;
            14'b11_001100011000: DATA = 12'b111101111110;
            14'b11_001100011001: DATA = 12'b111101111111;
            14'b11_001100011010: DATA = 12'b111110000000;
            14'b11_001100011011: DATA = 12'b111110000001;
            14'b11_001100011100: DATA = 12'b111110000011;
            14'b11_001100011101: DATA = 12'b111110000100;
            14'b11_001100011110: DATA = 12'b111110000101;
            14'b11_001100011111: DATA = 12'b111110000110;
            14'b11_001100100000: DATA = 12'b111110000111;
            14'b11_001100100001: DATA = 12'b111110001000;
            14'b11_001100100010: DATA = 12'b111110001001;
            14'b11_001100100011: DATA = 12'b111110001010;
            14'b11_001100100100: DATA = 12'b111110001011;
            14'b11_001100100101: DATA = 12'b111110001100;
            14'b11_001100100110: DATA = 12'b111110001101;
            14'b11_001100100111: DATA = 12'b111110001110;
            14'b11_001100101000: DATA = 12'b111110001111;
            14'b11_001100101001: DATA = 12'b111110010000;
            14'b11_001100101010: DATA = 12'b111110010001;
            14'b11_001100101011: DATA = 12'b111110010010;
            14'b11_001100101100: DATA = 12'b111110010011;
            14'b11_001100101101: DATA = 12'b111110010100;
            14'b11_001100101110: DATA = 12'b111110010101;
            14'b11_001100101111: DATA = 12'b111110010110;
            14'b11_001100110000: DATA = 12'b111110010111;
            14'b11_001100110001: DATA = 12'b111110011000;
            14'b11_001100110010: DATA = 12'b111110011001;
            14'b11_001100110011: DATA = 12'b111110011010;
            14'b11_001100110100: DATA = 12'b111110011011;
            14'b11_001100110101: DATA = 12'b111110011100;
            14'b11_001100110110: DATA = 12'b111110011101;
            14'b11_001100110111: DATA = 12'b111110011110;
            14'b11_001100111000: DATA = 12'b111110011111;
            14'b11_001100111001: DATA = 12'b111110100000;
            14'b11_001100111010: DATA = 12'b111110100001;
            14'b11_001100111011: DATA = 12'b111110100010;
            14'b11_001100111100: DATA = 12'b111110100011;
            14'b11_001100111101: DATA = 12'b111110100100;
            14'b11_001100111110: DATA = 12'b111110100101;
            14'b11_001100111111: DATA = 12'b111110100101;
            14'b11_001101000000: DATA = 12'b111110100110;
            14'b11_001101000001: DATA = 12'b111110100111;
            14'b11_001101000010: DATA = 12'b111110101000;
            14'b11_001101000011: DATA = 12'b111110101001;
            14'b11_001101000100: DATA = 12'b111110101010;
            14'b11_001101000101: DATA = 12'b111110101011;
            14'b11_001101000110: DATA = 12'b111110101100;
            14'b11_001101000111: DATA = 12'b111110101101;
            14'b11_001101001000: DATA = 12'b111110101110;
            14'b11_001101001001: DATA = 12'b111110101110;
            14'b11_001101001010: DATA = 12'b111110101111;
            14'b11_001101001011: DATA = 12'b111110110000;
            14'b11_001101001100: DATA = 12'b111110110001;
            14'b11_001101001101: DATA = 12'b111110110010;
            14'b11_001101001110: DATA = 12'b111110110011;
            14'b11_001101001111: DATA = 12'b111110110100;
            14'b11_001101010000: DATA = 12'b111110110100;
            14'b11_001101010001: DATA = 12'b111110110101;
            14'b11_001101010010: DATA = 12'b111110110110;
            14'b11_001101010011: DATA = 12'b111110110111;
            14'b11_001101010100: DATA = 12'b111110111000;
            14'b11_001101010101: DATA = 12'b111110111000;
            14'b11_001101010110: DATA = 12'b111110111001;
            14'b11_001101010111: DATA = 12'b111110111010;
            14'b11_001101011000: DATA = 12'b111110111011;
            14'b11_001101011001: DATA = 12'b111110111100;
            14'b11_001101011010: DATA = 12'b111110111100;
            14'b11_001101011011: DATA = 12'b111110111101;
            14'b11_001101011100: DATA = 12'b111110111110;
            14'b11_001101011101: DATA = 12'b111110111111;
            14'b11_001101011110: DATA = 12'b111111000000;
            14'b11_001101011111: DATA = 12'b111111000000;
            14'b11_001101100000: DATA = 12'b111111000001;
            14'b11_001101100001: DATA = 12'b111111000010;
            14'b11_001101100010: DATA = 12'b111111000011;
            14'b11_001101100011: DATA = 12'b111111000011;
            14'b11_001101100100: DATA = 12'b111111000100;
            14'b11_001101100101: DATA = 12'b111111000101;
            14'b11_001101100110: DATA = 12'b111111000110;
            14'b11_001101100111: DATA = 12'b111111000110;
            14'b11_001101101000: DATA = 12'b111111000111;
            14'b11_001101101001: DATA = 12'b111111001000;
            14'b11_001101101010: DATA = 12'b111111001001;
            14'b11_001101101011: DATA = 12'b111111001001;
            14'b11_001101101100: DATA = 12'b111111001010;
            14'b11_001101101101: DATA = 12'b111111001011;
            14'b11_001101101110: DATA = 12'b111111001011;
            14'b11_001101101111: DATA = 12'b111111001100;
            14'b11_001101110000: DATA = 12'b111111001101;
            14'b11_001101110001: DATA = 12'b111111001101;
            14'b11_001101110010: DATA = 12'b111111001110;
            14'b11_001101110011: DATA = 12'b111111001111;
            14'b11_001101110100: DATA = 12'b111111001111;
            14'b11_001101110101: DATA = 12'b111111010000;
            14'b11_001101110110: DATA = 12'b111111010001;
            14'b11_001101110111: DATA = 12'b111111010001;
            14'b11_001101111000: DATA = 12'b111111010010;
            14'b11_001101111001: DATA = 12'b111111010011;
            14'b11_001101111010: DATA = 12'b111111010011;
            14'b11_001101111011: DATA = 12'b111111010100;
            14'b11_001101111100: DATA = 12'b111111010101;
            14'b11_001101111101: DATA = 12'b111111010101;
            14'b11_001101111110: DATA = 12'b111111010110;
            14'b11_001101111111: DATA = 12'b111111010111;
            14'b11_001110000000: DATA = 12'b111111010111;
            14'b11_001110000001: DATA = 12'b111111011000;
            14'b11_001110000010: DATA = 12'b111111011000;
            14'b11_001110000011: DATA = 12'b111111011001;
            14'b11_001110000100: DATA = 12'b111111011010;
            14'b11_001110000101: DATA = 12'b111111011010;
            14'b11_001110000110: DATA = 12'b111111011011;
            14'b11_001110000111: DATA = 12'b111111011011;
            14'b11_001110001000: DATA = 12'b111111011100;
            14'b11_001110001001: DATA = 12'b111111011100;
            14'b11_001110001010: DATA = 12'b111111011101;
            14'b11_001110001011: DATA = 12'b111111011110;
            14'b11_001110001100: DATA = 12'b111111011110;
            14'b11_001110001101: DATA = 12'b111111011111;
            14'b11_001110001110: DATA = 12'b111111011111;
            14'b11_001110001111: DATA = 12'b111111100000;
            14'b11_001110010000: DATA = 12'b111111100000;
            14'b11_001110010001: DATA = 12'b111111100001;
            14'b11_001110010010: DATA = 12'b111111100001;
            14'b11_001110010011: DATA = 12'b111111100010;
            14'b11_001110010100: DATA = 12'b111111100010;
            14'b11_001110010101: DATA = 12'b111111100011;
            14'b11_001110010110: DATA = 12'b111111100011;
            14'b11_001110010111: DATA = 12'b111111100100;
            14'b11_001110011000: DATA = 12'b111111100101;
            14'b11_001110011001: DATA = 12'b111111100101;
            14'b11_001110011010: DATA = 12'b111111100101;
            14'b11_001110011011: DATA = 12'b111111100110;
            14'b11_001110011100: DATA = 12'b111111100110;
            14'b11_001110011101: DATA = 12'b111111100111;
            14'b11_001110011110: DATA = 12'b111111100111;
            14'b11_001110011111: DATA = 12'b111111101000;
            14'b11_001110100000: DATA = 12'b111111101000;
            14'b11_001110100001: DATA = 12'b111111101001;
            14'b11_001110100010: DATA = 12'b111111101001;
            14'b11_001110100011: DATA = 12'b111111101010;
            14'b11_001110100100: DATA = 12'b111111101010;
            14'b11_001110100101: DATA = 12'b111111101011;
            14'b11_001110100110: DATA = 12'b111111101011;
            14'b11_001110100111: DATA = 12'b111111101011;
            14'b11_001110101000: DATA = 12'b111111101100;
            14'b11_001110101001: DATA = 12'b111111101100;
            14'b11_001110101010: DATA = 12'b111111101101;
            14'b11_001110101011: DATA = 12'b111111101101;
            14'b11_001110101100: DATA = 12'b111111101110;
            14'b11_001110101101: DATA = 12'b111111101110;
            14'b11_001110101110: DATA = 12'b111111101110;
            14'b11_001110101111: DATA = 12'b111111101111;
            14'b11_001110110000: DATA = 12'b111111101111;
            14'b11_001110110001: DATA = 12'b111111101111;
            14'b11_001110110010: DATA = 12'b111111110000;
            14'b11_001110110011: DATA = 12'b111111110000;
            14'b11_001110110100: DATA = 12'b111111110001;
            14'b11_001110110101: DATA = 12'b111111110001;
            14'b11_001110110110: DATA = 12'b111111110001;
            14'b11_001110110111: DATA = 12'b111111110010;
            14'b11_001110111000: DATA = 12'b111111110010;
            14'b11_001110111001: DATA = 12'b111111110010;
            14'b11_001110111010: DATA = 12'b111111110011;
            14'b11_001110111011: DATA = 12'b111111110011;
            14'b11_001110111100: DATA = 12'b111111110011;
            14'b11_001110111101: DATA = 12'b111111110100;
            14'b11_001110111110: DATA = 12'b111111110100;
            14'b11_001110111111: DATA = 12'b111111110100;
            14'b11_001111000000: DATA = 12'b111111110101;
            14'b11_001111000001: DATA = 12'b111111110101;
            14'b11_001111000010: DATA = 12'b111111110101;
            14'b11_001111000011: DATA = 12'b111111110110;
            14'b11_001111000100: DATA = 12'b111111110110;
            14'b11_001111000101: DATA = 12'b111111110110;
            14'b11_001111000110: DATA = 12'b111111110110;
            14'b11_001111000111: DATA = 12'b111111110111;
            14'b11_001111001000: DATA = 12'b111111110111;
            14'b11_001111001001: DATA = 12'b111111110111;
            14'b11_001111001010: DATA = 12'b111111110111;
            14'b11_001111001011: DATA = 12'b111111111000;
            14'b11_001111001100: DATA = 12'b111111111000;
            14'b11_001111001101: DATA = 12'b111111111000;
            14'b11_001111001110: DATA = 12'b111111111000;
            14'b11_001111001111: DATA = 12'b111111111001;
            14'b11_001111010000: DATA = 12'b111111111001;
            14'b11_001111010001: DATA = 12'b111111111001;
            14'b11_001111010010: DATA = 12'b111111111001;
            14'b11_001111010011: DATA = 12'b111111111010;
            14'b11_001111010100: DATA = 12'b111111111010;
            14'b11_001111010101: DATA = 12'b111111111010;
            14'b11_001111010110: DATA = 12'b111111111010;
            14'b11_001111010111: DATA = 12'b111111111010;
            14'b11_001111011000: DATA = 12'b111111111011;
            14'b11_001111011001: DATA = 12'b111111111011;
            14'b11_001111011010: DATA = 12'b111111111011;
            14'b11_001111011011: DATA = 12'b111111111011;
            14'b11_001111011100: DATA = 12'b111111111011;
            14'b11_001111011101: DATA = 12'b111111111100;
            14'b11_001111011110: DATA = 12'b111111111100;
            14'b11_001111011111: DATA = 12'b111111111100;
            14'b11_001111100000: DATA = 12'b111111111100;
            14'b11_001111100001: DATA = 12'b111111111100;
            14'b11_001111100010: DATA = 12'b111111111100;
            14'b11_001111100011: DATA = 12'b111111111100;
            14'b11_001111100100: DATA = 12'b111111111101;
            14'b11_001111100101: DATA = 12'b111111111101;
            14'b11_001111100110: DATA = 12'b111111111101;
            14'b11_001111100111: DATA = 12'b111111111101;
            14'b11_001111101000: DATA = 12'b111111111101;
            14'b11_001111101001: DATA = 12'b111111111101;
            14'b11_001111101010: DATA = 12'b111111111101;
            14'b11_001111101011: DATA = 12'b111111111101;
            14'b11_001111101100: DATA = 12'b111111111110;
            14'b11_001111101101: DATA = 12'b111111111110;
            14'b11_001111101110: DATA = 12'b111111111110;
            14'b11_001111101111: DATA = 12'b111111111110;
            14'b11_001111110000: DATA = 12'b111111111110;
            14'b11_001111110001: DATA = 12'b111111111110;
            14'b11_001111110010: DATA = 12'b111111111110;
            14'b11_001111110011: DATA = 12'b111111111110;
            14'b11_001111110100: DATA = 12'b111111111110;
            14'b11_001111110101: DATA = 12'b111111111110;
            14'b11_001111110110: DATA = 12'b111111111110;
            14'b11_001111110111: DATA = 12'b111111111110;
            14'b11_001111111000: DATA = 12'b111111111110;
            14'b11_001111111001: DATA = 12'b111111111110;
            14'b11_001111111010: DATA = 12'b111111111110;
            14'b11_001111111011: DATA = 12'b111111111110;
            14'b11_001111111100: DATA = 12'b111111111110;
            14'b11_001111111101: DATA = 12'b111111111110;
            14'b11_001111111110: DATA = 12'b111111111110;
            14'b11_001111111111: DATA = 12'b111111111110;
            14'b11_010000000000: DATA = 12'b111111111111;
            14'b11_010000000001: DATA = 12'b111111111110;
            14'b11_010000000010: DATA = 12'b111111111110;
            14'b11_010000000011: DATA = 12'b111111111110;
            14'b11_010000000100: DATA = 12'b111111111110;
            14'b11_010000000101: DATA = 12'b111111111110;
            14'b11_010000000110: DATA = 12'b111111111110;
            14'b11_010000000111: DATA = 12'b111111111110;
            14'b11_010000001000: DATA = 12'b111111111110;
            14'b11_010000001001: DATA = 12'b111111111110;
            14'b11_010000001010: DATA = 12'b111111111110;
            14'b11_010000001011: DATA = 12'b111111111110;
            14'b11_010000001100: DATA = 12'b111111111110;
            14'b11_010000001101: DATA = 12'b111111111110;
            14'b11_010000001110: DATA = 12'b111111111110;
            14'b11_010000001111: DATA = 12'b111111111110;
            14'b11_010000010000: DATA = 12'b111111111110;
            14'b11_010000010001: DATA = 12'b111111111110;
            14'b11_010000010010: DATA = 12'b111111111110;
            14'b11_010000010011: DATA = 12'b111111111110;
            14'b11_010000010100: DATA = 12'b111111111110;
            14'b11_010000010101: DATA = 12'b111111111101;
            14'b11_010000010110: DATA = 12'b111111111101;
            14'b11_010000010111: DATA = 12'b111111111101;
            14'b11_010000011000: DATA = 12'b111111111101;
            14'b11_010000011001: DATA = 12'b111111111101;
            14'b11_010000011010: DATA = 12'b111111111101;
            14'b11_010000011011: DATA = 12'b111111111101;
            14'b11_010000011100: DATA = 12'b111111111101;
            14'b11_010000011101: DATA = 12'b111111111100;
            14'b11_010000011110: DATA = 12'b111111111100;
            14'b11_010000011111: DATA = 12'b111111111100;
            14'b11_010000100000: DATA = 12'b111111111100;
            14'b11_010000100001: DATA = 12'b111111111100;
            14'b11_010000100010: DATA = 12'b111111111100;
            14'b11_010000100011: DATA = 12'b111111111100;
            14'b11_010000100100: DATA = 12'b111111111011;
            14'b11_010000100101: DATA = 12'b111111111011;
            14'b11_010000100110: DATA = 12'b111111111011;
            14'b11_010000100111: DATA = 12'b111111111011;
            14'b11_010000101000: DATA = 12'b111111111011;
            14'b11_010000101001: DATA = 12'b111111111010;
            14'b11_010000101010: DATA = 12'b111111111010;
            14'b11_010000101011: DATA = 12'b111111111010;
            14'b11_010000101100: DATA = 12'b111111111010;
            14'b11_010000101101: DATA = 12'b111111111010;
            14'b11_010000101110: DATA = 12'b111111111001;
            14'b11_010000101111: DATA = 12'b111111111001;
            14'b11_010000110000: DATA = 12'b111111111001;
            14'b11_010000110001: DATA = 12'b111111111001;
            14'b11_010000110010: DATA = 12'b111111111000;
            14'b11_010000110011: DATA = 12'b111111111000;
            14'b11_010000110100: DATA = 12'b111111111000;
            14'b11_010000110101: DATA = 12'b111111111000;
            14'b11_010000110110: DATA = 12'b111111110111;
            14'b11_010000110111: DATA = 12'b111111110111;
            14'b11_010000111000: DATA = 12'b111111110111;
            14'b11_010000111001: DATA = 12'b111111110111;
            14'b11_010000111010: DATA = 12'b111111110110;
            14'b11_010000111011: DATA = 12'b111111110110;
            14'b11_010000111100: DATA = 12'b111111110110;
            14'b11_010000111101: DATA = 12'b111111110110;
            14'b11_010000111110: DATA = 12'b111111110101;
            14'b11_010000111111: DATA = 12'b111111110101;
            14'b11_010001000000: DATA = 12'b111111110101;
            14'b11_010001000001: DATA = 12'b111111110100;
            14'b11_010001000010: DATA = 12'b111111110100;
            14'b11_010001000011: DATA = 12'b111111110100;
            14'b11_010001000100: DATA = 12'b111111110011;
            14'b11_010001000101: DATA = 12'b111111110011;
            14'b11_010001000110: DATA = 12'b111111110011;
            14'b11_010001000111: DATA = 12'b111111110010;
            14'b11_010001001000: DATA = 12'b111111110010;
            14'b11_010001001001: DATA = 12'b111111110010;
            14'b11_010001001010: DATA = 12'b111111110001;
            14'b11_010001001011: DATA = 12'b111111110001;
            14'b11_010001001100: DATA = 12'b111111110001;
            14'b11_010001001101: DATA = 12'b111111110000;
            14'b11_010001001110: DATA = 12'b111111110000;
            14'b11_010001001111: DATA = 12'b111111101111;
            14'b11_010001010000: DATA = 12'b111111101111;
            14'b11_010001010001: DATA = 12'b111111101111;
            14'b11_010001010010: DATA = 12'b111111101110;
            14'b11_010001010011: DATA = 12'b111111101110;
            14'b11_010001010100: DATA = 12'b111111101110;
            14'b11_010001010101: DATA = 12'b111111101101;
            14'b11_010001010110: DATA = 12'b111111101101;
            14'b11_010001010111: DATA = 12'b111111101100;
            14'b11_010001011000: DATA = 12'b111111101100;
            14'b11_010001011001: DATA = 12'b111111101011;
            14'b11_010001011010: DATA = 12'b111111101011;
            14'b11_010001011011: DATA = 12'b111111101011;
            14'b11_010001011100: DATA = 12'b111111101010;
            14'b11_010001011101: DATA = 12'b111111101010;
            14'b11_010001011110: DATA = 12'b111111101001;
            14'b11_010001011111: DATA = 12'b111111101001;
            14'b11_010001100000: DATA = 12'b111111101000;
            14'b11_010001100001: DATA = 12'b111111101000;
            14'b11_010001100010: DATA = 12'b111111100111;
            14'b11_010001100011: DATA = 12'b111111100111;
            14'b11_010001100100: DATA = 12'b111111100110;
            14'b11_010001100101: DATA = 12'b111111100110;
            14'b11_010001100110: DATA = 12'b111111100101;
            14'b11_010001100111: DATA = 12'b111111100101;
            14'b11_010001101000: DATA = 12'b111111100101;
            14'b11_010001101001: DATA = 12'b111111100100;
            14'b11_010001101010: DATA = 12'b111111100011;
            14'b11_010001101011: DATA = 12'b111111100011;
            14'b11_010001101100: DATA = 12'b111111100010;
            14'b11_010001101101: DATA = 12'b111111100010;
            14'b11_010001101110: DATA = 12'b111111100001;
            14'b11_010001101111: DATA = 12'b111111100001;
            14'b11_010001110000: DATA = 12'b111111100000;
            14'b11_010001110001: DATA = 12'b111111100000;
            14'b11_010001110010: DATA = 12'b111111011111;
            14'b11_010001110011: DATA = 12'b111111011111;
            14'b11_010001110100: DATA = 12'b111111011110;
            14'b11_010001110101: DATA = 12'b111111011110;
            14'b11_010001110110: DATA = 12'b111111011101;
            14'b11_010001110111: DATA = 12'b111111011100;
            14'b11_010001111000: DATA = 12'b111111011100;
            14'b11_010001111001: DATA = 12'b111111011011;
            14'b11_010001111010: DATA = 12'b111111011011;
            14'b11_010001111011: DATA = 12'b111111011010;
            14'b11_010001111100: DATA = 12'b111111011010;
            14'b11_010001111101: DATA = 12'b111111011001;
            14'b11_010001111110: DATA = 12'b111111011000;
            14'b11_010001111111: DATA = 12'b111111011000;
            14'b11_010010000000: DATA = 12'b111111010111;
            14'b11_010010000001: DATA = 12'b111111010111;
            14'b11_010010000010: DATA = 12'b111111010110;
            14'b11_010010000011: DATA = 12'b111111010101;
            14'b11_010010000100: DATA = 12'b111111010101;
            14'b11_010010000101: DATA = 12'b111111010100;
            14'b11_010010000110: DATA = 12'b111111010011;
            14'b11_010010000111: DATA = 12'b111111010011;
            14'b11_010010001000: DATA = 12'b111111010010;
            14'b11_010010001001: DATA = 12'b111111010001;
            14'b11_010010001010: DATA = 12'b111111010001;
            14'b11_010010001011: DATA = 12'b111111010000;
            14'b11_010010001100: DATA = 12'b111111001111;
            14'b11_010010001101: DATA = 12'b111111001111;
            14'b11_010010001110: DATA = 12'b111111001110;
            14'b11_010010001111: DATA = 12'b111111001101;
            14'b11_010010010000: DATA = 12'b111111001101;
            14'b11_010010010001: DATA = 12'b111111001100;
            14'b11_010010010010: DATA = 12'b111111001011;
            14'b11_010010010011: DATA = 12'b111111001011;
            14'b11_010010010100: DATA = 12'b111111001010;
            14'b11_010010010101: DATA = 12'b111111001001;
            14'b11_010010010110: DATA = 12'b111111001001;
            14'b11_010010010111: DATA = 12'b111111001000;
            14'b11_010010011000: DATA = 12'b111111000111;
            14'b11_010010011001: DATA = 12'b111111000110;
            14'b11_010010011010: DATA = 12'b111111000110;
            14'b11_010010011011: DATA = 12'b111111000101;
            14'b11_010010011100: DATA = 12'b111111000100;
            14'b11_010010011101: DATA = 12'b111111000011;
            14'b11_010010011110: DATA = 12'b111111000011;
            14'b11_010010011111: DATA = 12'b111111000010;
            14'b11_010010100000: DATA = 12'b111111000001;
            14'b11_010010100001: DATA = 12'b111111000000;
            14'b11_010010100010: DATA = 12'b111111000000;
            14'b11_010010100011: DATA = 12'b111110111111;
            14'b11_010010100100: DATA = 12'b111110111110;
            14'b11_010010100101: DATA = 12'b111110111101;
            14'b11_010010100110: DATA = 12'b111110111100;
            14'b11_010010100111: DATA = 12'b111110111100;
            14'b11_010010101000: DATA = 12'b111110111011;
            14'b11_010010101001: DATA = 12'b111110111010;
            14'b11_010010101010: DATA = 12'b111110111001;
            14'b11_010010101011: DATA = 12'b111110111000;
            14'b11_010010101100: DATA = 12'b111110111000;
            14'b11_010010101101: DATA = 12'b111110110111;
            14'b11_010010101110: DATA = 12'b111110110110;
            14'b11_010010101111: DATA = 12'b111110110101;
            14'b11_010010110000: DATA = 12'b111110110100;
            14'b11_010010110001: DATA = 12'b111110110100;
            14'b11_010010110010: DATA = 12'b111110110011;
            14'b11_010010110011: DATA = 12'b111110110010;
            14'b11_010010110100: DATA = 12'b111110110001;
            14'b11_010010110101: DATA = 12'b111110110000;
            14'b11_010010110110: DATA = 12'b111110101111;
            14'b11_010010110111: DATA = 12'b111110101110;
            14'b11_010010111000: DATA = 12'b111110101110;
            14'b11_010010111001: DATA = 12'b111110101101;
            14'b11_010010111010: DATA = 12'b111110101100;
            14'b11_010010111011: DATA = 12'b111110101011;
            14'b11_010010111100: DATA = 12'b111110101010;
            14'b11_010010111101: DATA = 12'b111110101001;
            14'b11_010010111110: DATA = 12'b111110101000;
            14'b11_010010111111: DATA = 12'b111110100111;
            14'b11_010011000000: DATA = 12'b111110100110;
            14'b11_010011000001: DATA = 12'b111110100101;
            14'b11_010011000010: DATA = 12'b111110100101;
            14'b11_010011000011: DATA = 12'b111110100100;
            14'b11_010011000100: DATA = 12'b111110100011;
            14'b11_010011000101: DATA = 12'b111110100010;
            14'b11_010011000110: DATA = 12'b111110100001;
            14'b11_010011000111: DATA = 12'b111110100000;
            14'b11_010011001000: DATA = 12'b111110011111;
            14'b11_010011001001: DATA = 12'b111110011110;
            14'b11_010011001010: DATA = 12'b111110011101;
            14'b11_010011001011: DATA = 12'b111110011100;
            14'b11_010011001100: DATA = 12'b111110011011;
            14'b11_010011001101: DATA = 12'b111110011010;
            14'b11_010011001110: DATA = 12'b111110011001;
            14'b11_010011001111: DATA = 12'b111110011000;
            14'b11_010011010000: DATA = 12'b111110010111;
            14'b11_010011010001: DATA = 12'b111110010110;
            14'b11_010011010010: DATA = 12'b111110010101;
            14'b11_010011010011: DATA = 12'b111110010100;
            14'b11_010011010100: DATA = 12'b111110010011;
            14'b11_010011010101: DATA = 12'b111110010010;
            14'b11_010011010110: DATA = 12'b111110010001;
            14'b11_010011010111: DATA = 12'b111110010000;
            14'b11_010011011000: DATA = 12'b111110001111;
            14'b11_010011011001: DATA = 12'b111110001110;
            14'b11_010011011010: DATA = 12'b111110001101;
            14'b11_010011011011: DATA = 12'b111110001100;
            14'b11_010011011100: DATA = 12'b111110001011;
            14'b11_010011011101: DATA = 12'b111110001010;
            14'b11_010011011110: DATA = 12'b111110001001;
            14'b11_010011011111: DATA = 12'b111110001000;
            14'b11_010011100000: DATA = 12'b111110000111;
            14'b11_010011100001: DATA = 12'b111110000110;
            14'b11_010011100010: DATA = 12'b111110000101;
            14'b11_010011100011: DATA = 12'b111110000100;
            14'b11_010011100100: DATA = 12'b111110000011;
            14'b11_010011100101: DATA = 12'b111110000001;
            14'b11_010011100110: DATA = 12'b111110000000;
            14'b11_010011100111: DATA = 12'b111101111111;
            14'b11_010011101000: DATA = 12'b111101111110;
            14'b11_010011101001: DATA = 12'b111101111101;
            14'b11_010011101010: DATA = 12'b111101111100;
            14'b11_010011101011: DATA = 12'b111101111011;
            14'b11_010011101100: DATA = 12'b111101111010;
            14'b11_010011101101: DATA = 12'b111101111001;
            14'b11_010011101110: DATA = 12'b111101111000;
            14'b11_010011101111: DATA = 12'b111101110110;
            14'b11_010011110000: DATA = 12'b111101110101;
            14'b11_010011110001: DATA = 12'b111101110100;
            14'b11_010011110010: DATA = 12'b111101110011;
            14'b11_010011110011: DATA = 12'b111101110010;
            14'b11_010011110100: DATA = 12'b111101110001;
            14'b11_010011110101: DATA = 12'b111101110000;
            14'b11_010011110110: DATA = 12'b111101101110;
            14'b11_010011110111: DATA = 12'b111101101101;
            14'b11_010011111000: DATA = 12'b111101101100;
            14'b11_010011111001: DATA = 12'b111101101011;
            14'b11_010011111010: DATA = 12'b111101101010;
            14'b11_010011111011: DATA = 12'b111101101001;
            14'b11_010011111100: DATA = 12'b111101100111;
            14'b11_010011111101: DATA = 12'b111101100110;
            14'b11_010011111110: DATA = 12'b111101100101;
            14'b11_010011111111: DATA = 12'b111101100100;
            14'b11_010100000000: DATA = 12'b111101100011;
            14'b11_010100000001: DATA = 12'b111101100001;
            14'b11_010100000010: DATA = 12'b111101100000;
            14'b11_010100000011: DATA = 12'b111101011111;
            14'b11_010100000100: DATA = 12'b111101011110;
            14'b11_010100000101: DATA = 12'b111101011101;
            14'b11_010100000110: DATA = 12'b111101011011;
            14'b11_010100000111: DATA = 12'b111101011010;
            14'b11_010100001000: DATA = 12'b111101011001;
            14'b11_010100001001: DATA = 12'b111101011000;
            14'b11_010100001010: DATA = 12'b111101010110;
            14'b11_010100001011: DATA = 12'b111101010101;
            14'b11_010100001100: DATA = 12'b111101010100;
            14'b11_010100001101: DATA = 12'b111101010011;
            14'b11_010100001110: DATA = 12'b111101010001;
            14'b11_010100001111: DATA = 12'b111101010000;
            14'b11_010100010000: DATA = 12'b111101001111;
            14'b11_010100010001: DATA = 12'b111101001110;
            14'b11_010100010010: DATA = 12'b111101001100;
            14'b11_010100010011: DATA = 12'b111101001011;
            14'b11_010100010100: DATA = 12'b111101001010;
            14'b11_010100010101: DATA = 12'b111101001000;
            14'b11_010100010110: DATA = 12'b111101000111;
            14'b11_010100010111: DATA = 12'b111101000110;
            14'b11_010100011000: DATA = 12'b111101000101;
            14'b11_010100011001: DATA = 12'b111101000011;
            14'b11_010100011010: DATA = 12'b111101000010;
            14'b11_010100011011: DATA = 12'b111101000001;
            14'b11_010100011100: DATA = 12'b111100111111;
            14'b11_010100011101: DATA = 12'b111100111110;
            14'b11_010100011110: DATA = 12'b111100111101;
            14'b11_010100011111: DATA = 12'b111100111011;
            14'b11_010100100000: DATA = 12'b111100111010;
            14'b11_010100100001: DATA = 12'b111100111001;
            14'b11_010100100010: DATA = 12'b111100110111;
            14'b11_010100100011: DATA = 12'b111100110110;
            14'b11_010100100100: DATA = 12'b111100110101;
            14'b11_010100100101: DATA = 12'b111100110011;
            14'b11_010100100110: DATA = 12'b111100110010;
            14'b11_010100100111: DATA = 12'b111100110000;
            14'b11_010100101000: DATA = 12'b111100101111;
            14'b11_010100101001: DATA = 12'b111100101110;
            14'b11_010100101010: DATA = 12'b111100101100;
            14'b11_010100101011: DATA = 12'b111100101011;
            14'b11_010100101100: DATA = 12'b111100101010;
            14'b11_010100101101: DATA = 12'b111100101000;
            14'b11_010100101110: DATA = 12'b111100100111;
            14'b11_010100101111: DATA = 12'b111100100101;
            14'b11_010100110000: DATA = 12'b111100100100;
            14'b11_010100110001: DATA = 12'b111100100011;
            14'b11_010100110010: DATA = 12'b111100100001;
            14'b11_010100110011: DATA = 12'b111100100000;
            14'b11_010100110100: DATA = 12'b111100011110;
            14'b11_010100110101: DATA = 12'b111100011101;
            14'b11_010100110110: DATA = 12'b111100011011;
            14'b11_010100110111: DATA = 12'b111100011010;
            14'b11_010100111000: DATA = 12'b111100011000;
            14'b11_010100111001: DATA = 12'b111100010111;
            14'b11_010100111010: DATA = 12'b111100010110;
            14'b11_010100111011: DATA = 12'b111100010100;
            14'b11_010100111100: DATA = 12'b111100010011;
            14'b11_010100111101: DATA = 12'b111100010001;
            14'b11_010100111110: DATA = 12'b111100010000;
            14'b11_010100111111: DATA = 12'b111100001110;
            14'b11_010101000000: DATA = 12'b111100001101;
            14'b11_010101000001: DATA = 12'b111100001011;
            14'b11_010101000010: DATA = 12'b111100001010;
            14'b11_010101000011: DATA = 12'b111100001000;
            14'b11_010101000100: DATA = 12'b111100000111;
            14'b11_010101000101: DATA = 12'b111100000101;
            14'b11_010101000110: DATA = 12'b111100000100;
            14'b11_010101000111: DATA = 12'b111100000010;
            14'b11_010101001000: DATA = 12'b111100000001;
            14'b11_010101001001: DATA = 12'b111011111111;
            14'b11_010101001010: DATA = 12'b111011111110;
            14'b11_010101001011: DATA = 12'b111011111100;
            14'b11_010101001100: DATA = 12'b111011111011;
            14'b11_010101001101: DATA = 12'b111011111001;
            14'b11_010101001110: DATA = 12'b111011111000;
            14'b11_010101001111: DATA = 12'b111011110110;
            14'b11_010101010000: DATA = 12'b111011110101;
            14'b11_010101010001: DATA = 12'b111011110011;
            14'b11_010101010010: DATA = 12'b111011110001;
            14'b11_010101010011: DATA = 12'b111011110000;
            14'b11_010101010100: DATA = 12'b111011101110;
            14'b11_010101010101: DATA = 12'b111011101101;
            14'b11_010101010110: DATA = 12'b111011101011;
            14'b11_010101010111: DATA = 12'b111011101010;
            14'b11_010101011000: DATA = 12'b111011101000;
            14'b11_010101011001: DATA = 12'b111011100110;
            14'b11_010101011010: DATA = 12'b111011100101;
            14'b11_010101011011: DATA = 12'b111011100011;
            14'b11_010101011100: DATA = 12'b111011100010;
            14'b11_010101011101: DATA = 12'b111011100000;
            14'b11_010101011110: DATA = 12'b111011011110;
            14'b11_010101011111: DATA = 12'b111011011101;
            14'b11_010101100000: DATA = 12'b111011011011;
            14'b11_010101100001: DATA = 12'b111011011010;
            14'b11_010101100010: DATA = 12'b111011011000;
            14'b11_010101100011: DATA = 12'b111011010110;
            14'b11_010101100100: DATA = 12'b111011010101;
            14'b11_010101100101: DATA = 12'b111011010011;
            14'b11_010101100110: DATA = 12'b111011010010;
            14'b11_010101100111: DATA = 12'b111011010000;
            14'b11_010101101000: DATA = 12'b111011001110;
            14'b11_010101101001: DATA = 12'b111011001101;
            14'b11_010101101010: DATA = 12'b111011001011;
            14'b11_010101101011: DATA = 12'b111011001001;
            14'b11_010101101100: DATA = 12'b111011001000;
            14'b11_010101101101: DATA = 12'b111011000110;
            14'b11_010101101110: DATA = 12'b111011000100;
            14'b11_010101101111: DATA = 12'b111011000011;
            14'b11_010101110000: DATA = 12'b111011000001;
            14'b11_010101110001: DATA = 12'b111010111111;
            14'b11_010101110010: DATA = 12'b111010111110;
            14'b11_010101110011: DATA = 12'b111010111100;
            14'b11_010101110100: DATA = 12'b111010111010;
            14'b11_010101110101: DATA = 12'b111010111000;
            14'b11_010101110110: DATA = 12'b111010110111;
            14'b11_010101110111: DATA = 12'b111010110101;
            14'b11_010101111000: DATA = 12'b111010110011;
            14'b11_010101111001: DATA = 12'b111010110010;
            14'b11_010101111010: DATA = 12'b111010110000;
            14'b11_010101111011: DATA = 12'b111010101110;
            14'b11_010101111100: DATA = 12'b111010101100;
            14'b11_010101111101: DATA = 12'b111010101011;
            14'b11_010101111110: DATA = 12'b111010101001;
            14'b11_010101111111: DATA = 12'b111010100111;
            14'b11_010110000000: DATA = 12'b111010100110;
            14'b11_010110000001: DATA = 12'b111010100100;
            14'b11_010110000010: DATA = 12'b111010100010;
            14'b11_010110000011: DATA = 12'b111010100000;
            14'b11_010110000100: DATA = 12'b111010011111;
            14'b11_010110000101: DATA = 12'b111010011101;
            14'b11_010110000110: DATA = 12'b111010011011;
            14'b11_010110000111: DATA = 12'b111010011001;
            14'b11_010110001000: DATA = 12'b111010010111;
            14'b11_010110001001: DATA = 12'b111010010110;
            14'b11_010110001010: DATA = 12'b111010010100;
            14'b11_010110001011: DATA = 12'b111010010010;
            14'b11_010110001100: DATA = 12'b111010010000;
            14'b11_010110001101: DATA = 12'b111010001111;
            14'b11_010110001110: DATA = 12'b111010001101;
            14'b11_010110001111: DATA = 12'b111010001011;
            14'b11_010110010000: DATA = 12'b111010001001;
            14'b11_010110010001: DATA = 12'b111010000111;
            14'b11_010110010010: DATA = 12'b111010000101;
            14'b11_010110010011: DATA = 12'b111010000100;
            14'b11_010110010100: DATA = 12'b111010000010;
            14'b11_010110010101: DATA = 12'b111010000000;
            14'b11_010110010110: DATA = 12'b111001111110;
            14'b11_010110010111: DATA = 12'b111001111100;
            14'b11_010110011000: DATA = 12'b111001111011;
            14'b11_010110011001: DATA = 12'b111001111001;
            14'b11_010110011010: DATA = 12'b111001110111;
            14'b11_010110011011: DATA = 12'b111001110101;
            14'b11_010110011100: DATA = 12'b111001110011;
            14'b11_010110011101: DATA = 12'b111001110001;
            14'b11_010110011110: DATA = 12'b111001101111;
            14'b11_010110011111: DATA = 12'b111001101110;
            14'b11_010110100000: DATA = 12'b111001101100;
            14'b11_010110100001: DATA = 12'b111001101010;
            14'b11_010110100010: DATA = 12'b111001101000;
            14'b11_010110100011: DATA = 12'b111001100110;
            14'b11_010110100100: DATA = 12'b111001100100;
            14'b11_010110100101: DATA = 12'b111001100010;
            14'b11_010110100110: DATA = 12'b111001100000;
            14'b11_010110100111: DATA = 12'b111001011110;
            14'b11_010110101000: DATA = 12'b111001011101;
            14'b11_010110101001: DATA = 12'b111001011011;
            14'b11_010110101010: DATA = 12'b111001011001;
            14'b11_010110101011: DATA = 12'b111001010111;
            14'b11_010110101100: DATA = 12'b111001010101;
            14'b11_010110101101: DATA = 12'b111001010011;
            14'b11_010110101110: DATA = 12'b111001010001;
            14'b11_010110101111: DATA = 12'b111001001111;
            14'b11_010110110000: DATA = 12'b111001001101;
            14'b11_010110110001: DATA = 12'b111001001011;
            14'b11_010110110010: DATA = 12'b111001001001;
            14'b11_010110110011: DATA = 12'b111001000111;
            14'b11_010110110100: DATA = 12'b111001000101;
            14'b11_010110110101: DATA = 12'b111001000100;
            14'b11_010110110110: DATA = 12'b111001000010;
            14'b11_010110110111: DATA = 12'b111001000000;
            14'b11_010110111000: DATA = 12'b111000111110;
            14'b11_010110111001: DATA = 12'b111000111100;
            14'b11_010110111010: DATA = 12'b111000111010;
            14'b11_010110111011: DATA = 12'b111000111000;
            14'b11_010110111100: DATA = 12'b111000110110;
            14'b11_010110111101: DATA = 12'b111000110100;
            14'b11_010110111110: DATA = 12'b111000110010;
            14'b11_010110111111: DATA = 12'b111000110000;
            14'b11_010111000000: DATA = 12'b111000101110;
            14'b11_010111000001: DATA = 12'b111000101100;
            14'b11_010111000010: DATA = 12'b111000101010;
            14'b11_010111000011: DATA = 12'b111000101000;
            14'b11_010111000100: DATA = 12'b111000100110;
            14'b11_010111000101: DATA = 12'b111000100100;
            14'b11_010111000110: DATA = 12'b111000100010;
            14'b11_010111000111: DATA = 12'b111000100000;
            14'b11_010111001000: DATA = 12'b111000011110;
            14'b11_010111001001: DATA = 12'b111000011100;
            14'b11_010111001010: DATA = 12'b111000011010;
            14'b11_010111001011: DATA = 12'b111000011000;
            14'b11_010111001100: DATA = 12'b111000010110;
            14'b11_010111001101: DATA = 12'b111000010100;
            14'b11_010111001110: DATA = 12'b111000010010;
            14'b11_010111001111: DATA = 12'b111000010000;
            14'b11_010111010000: DATA = 12'b111000001110;
            14'b11_010111010001: DATA = 12'b111000001011;
            14'b11_010111010010: DATA = 12'b111000001001;
            14'b11_010111010011: DATA = 12'b111000000111;
            14'b11_010111010100: DATA = 12'b111000000101;
            14'b11_010111010101: DATA = 12'b111000000011;
            14'b11_010111010110: DATA = 12'b111000000001;
            14'b11_010111010111: DATA = 12'b110111111111;
            14'b11_010111011000: DATA = 12'b110111111101;
            14'b11_010111011001: DATA = 12'b110111111011;
            14'b11_010111011010: DATA = 12'b110111111001;
            14'b11_010111011011: DATA = 12'b110111110111;
            14'b11_010111011100: DATA = 12'b110111110101;
            14'b11_010111011101: DATA = 12'b110111110011;
            14'b11_010111011110: DATA = 12'b110111110000;
            14'b11_010111011111: DATA = 12'b110111101110;
            14'b11_010111100000: DATA = 12'b110111101100;
            14'b11_010111100001: DATA = 12'b110111101010;
            14'b11_010111100010: DATA = 12'b110111101000;
            14'b11_010111100011: DATA = 12'b110111100110;
            14'b11_010111100100: DATA = 12'b110111100100;
            14'b11_010111100101: DATA = 12'b110111100010;
            14'b11_010111100110: DATA = 12'b110111100000;
            14'b11_010111100111: DATA = 12'b110111011101;
            14'b11_010111101000: DATA = 12'b110111011011;
            14'b11_010111101001: DATA = 12'b110111011001;
            14'b11_010111101010: DATA = 12'b110111010111;
            14'b11_010111101011: DATA = 12'b110111010101;
            14'b11_010111101100: DATA = 12'b110111010011;
            14'b11_010111101101: DATA = 12'b110111010001;
            14'b11_010111101110: DATA = 12'b110111001110;
            14'b11_010111101111: DATA = 12'b110111001100;
            14'b11_010111110000: DATA = 12'b110111001010;
            14'b11_010111110001: DATA = 12'b110111001000;
            14'b11_010111110010: DATA = 12'b110111000110;
            14'b11_010111110011: DATA = 12'b110111000100;
            14'b11_010111110100: DATA = 12'b110111000001;
            14'b11_010111110101: DATA = 12'b110110111111;
            14'b11_010111110110: DATA = 12'b110110111101;
            14'b11_010111110111: DATA = 12'b110110111011;
            14'b11_010111111000: DATA = 12'b110110111001;
            14'b11_010111111001: DATA = 12'b110110110110;
            14'b11_010111111010: DATA = 12'b110110110100;
            14'b11_010111111011: DATA = 12'b110110110010;
            14'b11_010111111100: DATA = 12'b110110110000;
            14'b11_010111111101: DATA = 12'b110110101110;
            14'b11_010111111110: DATA = 12'b110110101011;
            14'b11_010111111111: DATA = 12'b110110101001;
            14'b11_011000000000: DATA = 12'b110110100111;
            14'b11_011000000001: DATA = 12'b110110100101;
            14'b11_011000000010: DATA = 12'b110110100011;
            14'b11_011000000011: DATA = 12'b110110100000;
            14'b11_011000000100: DATA = 12'b110110011110;
            14'b11_011000000101: DATA = 12'b110110011100;
            14'b11_011000000110: DATA = 12'b110110011010;
            14'b11_011000000111: DATA = 12'b110110010111;
            14'b11_011000001000: DATA = 12'b110110010101;
            14'b11_011000001001: DATA = 12'b110110010011;
            14'b11_011000001010: DATA = 12'b110110010001;
            14'b11_011000001011: DATA = 12'b110110001110;
            14'b11_011000001100: DATA = 12'b110110001100;
            14'b11_011000001101: DATA = 12'b110110001010;
            14'b11_011000001110: DATA = 12'b110110001000;
            14'b11_011000001111: DATA = 12'b110110000101;
            14'b11_011000010000: DATA = 12'b110110000011;
            14'b11_011000010001: DATA = 12'b110110000001;
            14'b11_011000010010: DATA = 12'b110101111110;
            14'b11_011000010011: DATA = 12'b110101111100;
            14'b11_011000010100: DATA = 12'b110101111010;
            14'b11_011000010101: DATA = 12'b110101111000;
            14'b11_011000010110: DATA = 12'b110101110101;
            14'b11_011000010111: DATA = 12'b110101110011;
            14'b11_011000011000: DATA = 12'b110101110001;
            14'b11_011000011001: DATA = 12'b110101101110;
            14'b11_011000011010: DATA = 12'b110101101100;
            14'b11_011000011011: DATA = 12'b110101101010;
            14'b11_011000011100: DATA = 12'b110101100111;
            14'b11_011000011101: DATA = 12'b110101100101;
            14'b11_011000011110: DATA = 12'b110101100011;
            14'b11_011000011111: DATA = 12'b110101100001;
            14'b11_011000100000: DATA = 12'b110101011110;
            14'b11_011000100001: DATA = 12'b110101011100;
            14'b11_011000100010: DATA = 12'b110101011010;
            14'b11_011000100011: DATA = 12'b110101010111;
            14'b11_011000100100: DATA = 12'b110101010101;
            14'b11_011000100101: DATA = 12'b110101010011;
            14'b11_011000100110: DATA = 12'b110101010000;
            14'b11_011000100111: DATA = 12'b110101001110;
            14'b11_011000101000: DATA = 12'b110101001011;
            14'b11_011000101001: DATA = 12'b110101001001;
            14'b11_011000101010: DATA = 12'b110101000111;
            14'b11_011000101011: DATA = 12'b110101000100;
            14'b11_011000101100: DATA = 12'b110101000010;
            14'b11_011000101101: DATA = 12'b110101000000;
            14'b11_011000101110: DATA = 12'b110100111101;
            14'b11_011000101111: DATA = 12'b110100111011;
            14'b11_011000110000: DATA = 12'b110100111001;
            14'b11_011000110001: DATA = 12'b110100110110;
            14'b11_011000110010: DATA = 12'b110100110100;
            14'b11_011000110011: DATA = 12'b110100110001;
            14'b11_011000110100: DATA = 12'b110100101111;
            14'b11_011000110101: DATA = 12'b110100101101;
            14'b11_011000110110: DATA = 12'b110100101010;
            14'b11_011000110111: DATA = 12'b110100101000;
            14'b11_011000111000: DATA = 12'b110100100101;
            14'b11_011000111001: DATA = 12'b110100100011;
            14'b11_011000111010: DATA = 12'b110100100001;
            14'b11_011000111011: DATA = 12'b110100011110;
            14'b11_011000111100: DATA = 12'b110100011100;
            14'b11_011000111101: DATA = 12'b110100011001;
            14'b11_011000111110: DATA = 12'b110100010111;
            14'b11_011000111111: DATA = 12'b110100010101;
            14'b11_011001000000: DATA = 12'b110100010010;
            14'b11_011001000001: DATA = 12'b110100010000;
            14'b11_011001000010: DATA = 12'b110100001101;
            14'b11_011001000011: DATA = 12'b110100001011;
            14'b11_011001000100: DATA = 12'b110100001000;
            14'b11_011001000101: DATA = 12'b110100000110;
            14'b11_011001000110: DATA = 12'b110100000011;
            14'b11_011001000111: DATA = 12'b110100000001;
            14'b11_011001001000: DATA = 12'b110011111111;
            14'b11_011001001001: DATA = 12'b110011111100;
            14'b11_011001001010: DATA = 12'b110011111010;
            14'b11_011001001011: DATA = 12'b110011110111;
            14'b11_011001001100: DATA = 12'b110011110101;
            14'b11_011001001101: DATA = 12'b110011110010;
            14'b11_011001001110: DATA = 12'b110011110000;
            14'b11_011001001111: DATA = 12'b110011101101;
            14'b11_011001010000: DATA = 12'b110011101011;
            14'b11_011001010001: DATA = 12'b110011101000;
            14'b11_011001010010: DATA = 12'b110011100110;
            14'b11_011001010011: DATA = 12'b110011100011;
            14'b11_011001010100: DATA = 12'b110011100001;
            14'b11_011001010101: DATA = 12'b110011011110;
            14'b11_011001010110: DATA = 12'b110011011100;
            14'b11_011001010111: DATA = 12'b110011011001;
            14'b11_011001011000: DATA = 12'b110011010111;
            14'b11_011001011001: DATA = 12'b110011010100;
            14'b11_011001011010: DATA = 12'b110011010010;
            14'b11_011001011011: DATA = 12'b110011001111;
            14'b11_011001011100: DATA = 12'b110011001101;
            14'b11_011001011101: DATA = 12'b110011001010;
            14'b11_011001011110: DATA = 12'b110011001000;
            14'b11_011001011111: DATA = 12'b110011000101;
            14'b11_011001100000: DATA = 12'b110011000011;
            14'b11_011001100001: DATA = 12'b110011000000;
            14'b11_011001100010: DATA = 12'b110010111110;
            14'b11_011001100011: DATA = 12'b110010111011;
            14'b11_011001100100: DATA = 12'b110010111001;
            14'b11_011001100101: DATA = 12'b110010110110;
            14'b11_011001100110: DATA = 12'b110010110100;
            14'b11_011001100111: DATA = 12'b110010110001;
            14'b11_011001101000: DATA = 12'b110010101111;
            14'b11_011001101001: DATA = 12'b110010101100;
            14'b11_011001101010: DATA = 12'b110010101010;
            14'b11_011001101011: DATA = 12'b110010100111;
            14'b11_011001101100: DATA = 12'b110010100100;
            14'b11_011001101101: DATA = 12'b110010100010;
            14'b11_011001101110: DATA = 12'b110010011111;
            14'b11_011001101111: DATA = 12'b110010011101;
            14'b11_011001110000: DATA = 12'b110010011010;
            14'b11_011001110001: DATA = 12'b110010011000;
            14'b11_011001110010: DATA = 12'b110010010101;
            14'b11_011001110011: DATA = 12'b110010010010;
            14'b11_011001110100: DATA = 12'b110010010000;
            14'b11_011001110101: DATA = 12'b110010001101;
            14'b11_011001110110: DATA = 12'b110010001011;
            14'b11_011001110111: DATA = 12'b110010001000;
            14'b11_011001111000: DATA = 12'b110010000110;
            14'b11_011001111001: DATA = 12'b110010000011;
            14'b11_011001111010: DATA = 12'b110010000000;
            14'b11_011001111011: DATA = 12'b110001111110;
            14'b11_011001111100: DATA = 12'b110001111011;
            14'b11_011001111101: DATA = 12'b110001111001;
            14'b11_011001111110: DATA = 12'b110001110110;
            14'b11_011001111111: DATA = 12'b110001110011;
            14'b11_011010000000: DATA = 12'b110001110001;
            14'b11_011010000001: DATA = 12'b110001101110;
            14'b11_011010000010: DATA = 12'b110001101100;
            14'b11_011010000011: DATA = 12'b110001101001;
            14'b11_011010000100: DATA = 12'b110001100110;
            14'b11_011010000101: DATA = 12'b110001100100;
            14'b11_011010000110: DATA = 12'b110001100001;
            14'b11_011010000111: DATA = 12'b110001011110;
            14'b11_011010001000: DATA = 12'b110001011100;
            14'b11_011010001001: DATA = 12'b110001011001;
            14'b11_011010001010: DATA = 12'b110001010111;
            14'b11_011010001011: DATA = 12'b110001010100;
            14'b11_011010001100: DATA = 12'b110001010001;
            14'b11_011010001101: DATA = 12'b110001001111;
            14'b11_011010001110: DATA = 12'b110001001100;
            14'b11_011010001111: DATA = 12'b110001001001;
            14'b11_011010010000: DATA = 12'b110001000111;
            14'b11_011010010001: DATA = 12'b110001000100;
            14'b11_011010010010: DATA = 12'b110001000001;
            14'b11_011010010011: DATA = 12'b110000111111;
            14'b11_011010010100: DATA = 12'b110000111100;
            14'b11_011010010101: DATA = 12'b110000111001;
            14'b11_011010010110: DATA = 12'b110000110111;
            14'b11_011010010111: DATA = 12'b110000110100;
            14'b11_011010011000: DATA = 12'b110000110001;
            14'b11_011010011001: DATA = 12'b110000101111;
            14'b11_011010011010: DATA = 12'b110000101100;
            14'b11_011010011011: DATA = 12'b110000101001;
            14'b11_011010011100: DATA = 12'b110000100111;
            14'b11_011010011101: DATA = 12'b110000100100;
            14'b11_011010011110: DATA = 12'b110000100001;
            14'b11_011010011111: DATA = 12'b110000011111;
            14'b11_011010100000: DATA = 12'b110000011100;
            14'b11_011010100001: DATA = 12'b110000011001;
            14'b11_011010100010: DATA = 12'b110000010110;
            14'b11_011010100011: DATA = 12'b110000010100;
            14'b11_011010100100: DATA = 12'b110000010001;
            14'b11_011010100101: DATA = 12'b110000001110;
            14'b11_011010100110: DATA = 12'b110000001100;
            14'b11_011010100111: DATA = 12'b110000001001;
            14'b11_011010101000: DATA = 12'b110000000110;
            14'b11_011010101001: DATA = 12'b110000000100;
            14'b11_011010101010: DATA = 12'b110000000001;
            14'b11_011010101011: DATA = 12'b101111111110;
            14'b11_011010101100: DATA = 12'b101111111011;
            14'b11_011010101101: DATA = 12'b101111111001;
            14'b11_011010101110: DATA = 12'b101111110110;
            14'b11_011010101111: DATA = 12'b101111110011;
            14'b11_011010110000: DATA = 12'b101111110000;
            14'b11_011010110001: DATA = 12'b101111101110;
            14'b11_011010110010: DATA = 12'b101111101011;
            14'b11_011010110011: DATA = 12'b101111101000;
            14'b11_011010110100: DATA = 12'b101111100110;
            14'b11_011010110101: DATA = 12'b101111100011;
            14'b11_011010110110: DATA = 12'b101111100000;
            14'b11_011010110111: DATA = 12'b101111011101;
            14'b11_011010111000: DATA = 12'b101111011011;
            14'b11_011010111001: DATA = 12'b101111011000;
            14'b11_011010111010: DATA = 12'b101111010101;
            14'b11_011010111011: DATA = 12'b101111010010;
            14'b11_011010111100: DATA = 12'b101111010000;
            14'b11_011010111101: DATA = 12'b101111001101;
            14'b11_011010111110: DATA = 12'b101111001010;
            14'b11_011010111111: DATA = 12'b101111000111;
            14'b11_011011000000: DATA = 12'b101111000100;
            14'b11_011011000001: DATA = 12'b101111000010;
            14'b11_011011000010: DATA = 12'b101110111111;
            14'b11_011011000011: DATA = 12'b101110111100;
            14'b11_011011000100: DATA = 12'b101110111001;
            14'b11_011011000101: DATA = 12'b101110110111;
            14'b11_011011000110: DATA = 12'b101110110100;
            14'b11_011011000111: DATA = 12'b101110110001;
            14'b11_011011001000: DATA = 12'b101110101110;
            14'b11_011011001001: DATA = 12'b101110101011;
            14'b11_011011001010: DATA = 12'b101110101001;
            14'b11_011011001011: DATA = 12'b101110100110;
            14'b11_011011001100: DATA = 12'b101110100011;
            14'b11_011011001101: DATA = 12'b101110100000;
            14'b11_011011001110: DATA = 12'b101110011101;
            14'b11_011011001111: DATA = 12'b101110011011;
            14'b11_011011010000: DATA = 12'b101110011000;
            14'b11_011011010001: DATA = 12'b101110010101;
            14'b11_011011010010: DATA = 12'b101110010010;
            14'b11_011011010011: DATA = 12'b101110001111;
            14'b11_011011010100: DATA = 12'b101110001101;
            14'b11_011011010101: DATA = 12'b101110001010;
            14'b11_011011010110: DATA = 12'b101110000111;
            14'b11_011011010111: DATA = 12'b101110000100;
            14'b11_011011011000: DATA = 12'b101110000001;
            14'b11_011011011001: DATA = 12'b101101111111;
            14'b11_011011011010: DATA = 12'b101101111100;
            14'b11_011011011011: DATA = 12'b101101111001;
            14'b11_011011011100: DATA = 12'b101101110110;
            14'b11_011011011101: DATA = 12'b101101110011;
            14'b11_011011011110: DATA = 12'b101101110000;
            14'b11_011011011111: DATA = 12'b101101101110;
            14'b11_011011100000: DATA = 12'b101101101011;
            14'b11_011011100001: DATA = 12'b101101101000;
            14'b11_011011100010: DATA = 12'b101101100101;
            14'b11_011011100011: DATA = 12'b101101100010;
            14'b11_011011100100: DATA = 12'b101101011111;
            14'b11_011011100101: DATA = 12'b101101011100;
            14'b11_011011100110: DATA = 12'b101101011010;
            14'b11_011011100111: DATA = 12'b101101010111;
            14'b11_011011101000: DATA = 12'b101101010100;
            14'b11_011011101001: DATA = 12'b101101010001;
            14'b11_011011101010: DATA = 12'b101101001110;
            14'b11_011011101011: DATA = 12'b101101001011;
            14'b11_011011101100: DATA = 12'b101101001000;
            14'b11_011011101101: DATA = 12'b101101000110;
            14'b11_011011101110: DATA = 12'b101101000011;
            14'b11_011011101111: DATA = 12'b101101000000;
            14'b11_011011110000: DATA = 12'b101100111101;
            14'b11_011011110001: DATA = 12'b101100111010;
            14'b11_011011110010: DATA = 12'b101100110111;
            14'b11_011011110011: DATA = 12'b101100110100;
            14'b11_011011110100: DATA = 12'b101100110010;
            14'b11_011011110101: DATA = 12'b101100101111;
            14'b11_011011110110: DATA = 12'b101100101100;
            14'b11_011011110111: DATA = 12'b101100101001;
            14'b11_011011111000: DATA = 12'b101100100110;
            14'b11_011011111001: DATA = 12'b101100100011;
            14'b11_011011111010: DATA = 12'b101100100000;
            14'b11_011011111011: DATA = 12'b101100011101;
            14'b11_011011111100: DATA = 12'b101100011010;
            14'b11_011011111101: DATA = 12'b101100011000;
            14'b11_011011111110: DATA = 12'b101100010101;
            14'b11_011011111111: DATA = 12'b101100010010;
            14'b11_011100000000: DATA = 12'b101100001111;
            14'b11_011100000001: DATA = 12'b101100001100;
            14'b11_011100000010: DATA = 12'b101100001001;
            14'b11_011100000011: DATA = 12'b101100000110;
            14'b11_011100000100: DATA = 12'b101100000011;
            14'b11_011100000101: DATA = 12'b101100000000;
            14'b11_011100000110: DATA = 12'b101011111101;
            14'b11_011100000111: DATA = 12'b101011111011;
            14'b11_011100001000: DATA = 12'b101011111000;
            14'b11_011100001001: DATA = 12'b101011110101;
            14'b11_011100001010: DATA = 12'b101011110010;
            14'b11_011100001011: DATA = 12'b101011101111;
            14'b11_011100001100: DATA = 12'b101011101100;
            14'b11_011100001101: DATA = 12'b101011101001;
            14'b11_011100001110: DATA = 12'b101011100110;
            14'b11_011100001111: DATA = 12'b101011100011;
            14'b11_011100010000: DATA = 12'b101011100000;
            14'b11_011100010001: DATA = 12'b101011011101;
            14'b11_011100010010: DATA = 12'b101011011010;
            14'b11_011100010011: DATA = 12'b101011010111;
            14'b11_011100010100: DATA = 12'b101011010100;
            14'b11_011100010101: DATA = 12'b101011010010;
            14'b11_011100010110: DATA = 12'b101011001111;
            14'b11_011100010111: DATA = 12'b101011001100;
            14'b11_011100011000: DATA = 12'b101011001001;
            14'b11_011100011001: DATA = 12'b101011000110;
            14'b11_011100011010: DATA = 12'b101011000011;
            14'b11_011100011011: DATA = 12'b101011000000;
            14'b11_011100011100: DATA = 12'b101010111101;
            14'b11_011100011101: DATA = 12'b101010111010;
            14'b11_011100011110: DATA = 12'b101010110111;
            14'b11_011100011111: DATA = 12'b101010110100;
            14'b11_011100100000: DATA = 12'b101010110001;
            14'b11_011100100001: DATA = 12'b101010101110;
            14'b11_011100100010: DATA = 12'b101010101011;
            14'b11_011100100011: DATA = 12'b101010101000;
            14'b11_011100100100: DATA = 12'b101010100101;
            14'b11_011100100101: DATA = 12'b101010100010;
            14'b11_011100100110: DATA = 12'b101010011111;
            14'b11_011100100111: DATA = 12'b101010011100;
            14'b11_011100101000: DATA = 12'b101010011001;
            14'b11_011100101001: DATA = 12'b101010010110;
            14'b11_011100101010: DATA = 12'b101010010011;
            14'b11_011100101011: DATA = 12'b101010010000;
            14'b11_011100101100: DATA = 12'b101010001110;
            14'b11_011100101101: DATA = 12'b101010001011;
            14'b11_011100101110: DATA = 12'b101010001000;
            14'b11_011100101111: DATA = 12'b101010000101;
            14'b11_011100110000: DATA = 12'b101010000010;
            14'b11_011100110001: DATA = 12'b101001111111;
            14'b11_011100110010: DATA = 12'b101001111100;
            14'b11_011100110011: DATA = 12'b101001111001;
            14'b11_011100110100: DATA = 12'b101001110110;
            14'b11_011100110101: DATA = 12'b101001110011;
            14'b11_011100110110: DATA = 12'b101001110000;
            14'b11_011100110111: DATA = 12'b101001101101;
            14'b11_011100111000: DATA = 12'b101001101010;
            14'b11_011100111001: DATA = 12'b101001100111;
            14'b11_011100111010: DATA = 12'b101001100100;
            14'b11_011100111011: DATA = 12'b101001100001;
            14'b11_011100111100: DATA = 12'b101001011110;
            14'b11_011100111101: DATA = 12'b101001011011;
            14'b11_011100111110: DATA = 12'b101001011000;
            14'b11_011100111111: DATA = 12'b101001010101;
            14'b11_011101000000: DATA = 12'b101001010010;
            14'b11_011101000001: DATA = 12'b101001001111;
            14'b11_011101000010: DATA = 12'b101001001100;
            14'b11_011101000011: DATA = 12'b101001001001;
            14'b11_011101000100: DATA = 12'b101001000110;
            14'b11_011101000101: DATA = 12'b101001000011;
            14'b11_011101000110: DATA = 12'b101001000000;
            14'b11_011101000111: DATA = 12'b101000111101;
            14'b11_011101001000: DATA = 12'b101000111010;
            14'b11_011101001001: DATA = 12'b101000110111;
            14'b11_011101001010: DATA = 12'b101000110100;
            14'b11_011101001011: DATA = 12'b101000110001;
            14'b11_011101001100: DATA = 12'b101000101110;
            14'b11_011101001101: DATA = 12'b101000101011;
            14'b11_011101001110: DATA = 12'b101000101000;
            14'b11_011101001111: DATA = 12'b101000100100;
            14'b11_011101010000: DATA = 12'b101000100001;
            14'b11_011101010001: DATA = 12'b101000011110;
            14'b11_011101010010: DATA = 12'b101000011011;
            14'b11_011101010011: DATA = 12'b101000011000;
            14'b11_011101010100: DATA = 12'b101000010101;
            14'b11_011101010101: DATA = 12'b101000010010;
            14'b11_011101010110: DATA = 12'b101000001111;
            14'b11_011101010111: DATA = 12'b101000001100;
            14'b11_011101011000: DATA = 12'b101000001001;
            14'b11_011101011001: DATA = 12'b101000000110;
            14'b11_011101011010: DATA = 12'b101000000011;
            14'b11_011101011011: DATA = 12'b101000000000;
            14'b11_011101011100: DATA = 12'b100111111101;
            14'b11_011101011101: DATA = 12'b100111111010;
            14'b11_011101011110: DATA = 12'b100111110111;
            14'b11_011101011111: DATA = 12'b100111110100;
            14'b11_011101100000: DATA = 12'b100111110001;
            14'b11_011101100001: DATA = 12'b100111101110;
            14'b11_011101100010: DATA = 12'b100111101011;
            14'b11_011101100011: DATA = 12'b100111101000;
            14'b11_011101100100: DATA = 12'b100111100101;
            14'b11_011101100101: DATA = 12'b100111100010;
            14'b11_011101100110: DATA = 12'b100111011111;
            14'b11_011101100111: DATA = 12'b100111011100;
            14'b11_011101101000: DATA = 12'b100111011000;
            14'b11_011101101001: DATA = 12'b100111010101;
            14'b11_011101101010: DATA = 12'b100111010010;
            14'b11_011101101011: DATA = 12'b100111001111;
            14'b11_011101101100: DATA = 12'b100111001100;
            14'b11_011101101101: DATA = 12'b100111001001;
            14'b11_011101101110: DATA = 12'b100111000110;
            14'b11_011101101111: DATA = 12'b100111000011;
            14'b11_011101110000: DATA = 12'b100111000000;
            14'b11_011101110001: DATA = 12'b100110111101;
            14'b11_011101110010: DATA = 12'b100110111010;
            14'b11_011101110011: DATA = 12'b100110110111;
            14'b11_011101110100: DATA = 12'b100110110100;
            14'b11_011101110101: DATA = 12'b100110110001;
            14'b11_011101110110: DATA = 12'b100110101110;
            14'b11_011101110111: DATA = 12'b100110101011;
            14'b11_011101111000: DATA = 12'b100110100111;
            14'b11_011101111001: DATA = 12'b100110100100;
            14'b11_011101111010: DATA = 12'b100110100001;
            14'b11_011101111011: DATA = 12'b100110011110;
            14'b11_011101111100: DATA = 12'b100110011011;
            14'b11_011101111101: DATA = 12'b100110011000;
            14'b11_011101111110: DATA = 12'b100110010101;
            14'b11_011101111111: DATA = 12'b100110010010;
            14'b11_011110000000: DATA = 12'b100110001111;
            14'b11_011110000001: DATA = 12'b100110001100;
            14'b11_011110000010: DATA = 12'b100110001001;
            14'b11_011110000011: DATA = 12'b100110000110;
            14'b11_011110000100: DATA = 12'b100110000011;
            14'b11_011110000101: DATA = 12'b100101111111;
            14'b11_011110000110: DATA = 12'b100101111100;
            14'b11_011110000111: DATA = 12'b100101111001;
            14'b11_011110001000: DATA = 12'b100101110110;
            14'b11_011110001001: DATA = 12'b100101110011;
            14'b11_011110001010: DATA = 12'b100101110000;
            14'b11_011110001011: DATA = 12'b100101101101;
            14'b11_011110001100: DATA = 12'b100101101010;
            14'b11_011110001101: DATA = 12'b100101100111;
            14'b11_011110001110: DATA = 12'b100101100100;
            14'b11_011110001111: DATA = 12'b100101100001;
            14'b11_011110010000: DATA = 12'b100101011101;
            14'b11_011110010001: DATA = 12'b100101011010;
            14'b11_011110010010: DATA = 12'b100101010111;
            14'b11_011110010011: DATA = 12'b100101010100;
            14'b11_011110010100: DATA = 12'b100101010001;
            14'b11_011110010101: DATA = 12'b100101001110;
            14'b11_011110010110: DATA = 12'b100101001011;
            14'b11_011110010111: DATA = 12'b100101001000;
            14'b11_011110011000: DATA = 12'b100101000101;
            14'b11_011110011001: DATA = 12'b100101000010;
            14'b11_011110011010: DATA = 12'b100100111110;
            14'b11_011110011011: DATA = 12'b100100111011;
            14'b11_011110011100: DATA = 12'b100100111000;
            14'b11_011110011101: DATA = 12'b100100110101;
            14'b11_011110011110: DATA = 12'b100100110010;
            14'b11_011110011111: DATA = 12'b100100101111;
            14'b11_011110100000: DATA = 12'b100100101100;
            14'b11_011110100001: DATA = 12'b100100101001;
            14'b11_011110100010: DATA = 12'b100100100110;
            14'b11_011110100011: DATA = 12'b100100100011;
            14'b11_011110100100: DATA = 12'b100100011111;
            14'b11_011110100101: DATA = 12'b100100011100;
            14'b11_011110100110: DATA = 12'b100100011001;
            14'b11_011110100111: DATA = 12'b100100010110;
            14'b11_011110101000: DATA = 12'b100100010011;
            14'b11_011110101001: DATA = 12'b100100010000;
            14'b11_011110101010: DATA = 12'b100100001101;
            14'b11_011110101011: DATA = 12'b100100001010;
            14'b11_011110101100: DATA = 12'b100100000111;
            14'b11_011110101101: DATA = 12'b100100000011;
            14'b11_011110101110: DATA = 12'b100100000000;
            14'b11_011110101111: DATA = 12'b100011111101;
            14'b11_011110110000: DATA = 12'b100011111010;
            14'b11_011110110001: DATA = 12'b100011110111;
            14'b11_011110110010: DATA = 12'b100011110100;
            14'b11_011110110011: DATA = 12'b100011110001;
            14'b11_011110110100: DATA = 12'b100011101110;
            14'b11_011110110101: DATA = 12'b100011101010;
            14'b11_011110110110: DATA = 12'b100011100111;
            14'b11_011110110111: DATA = 12'b100011100100;
            14'b11_011110111000: DATA = 12'b100011100001;
            14'b11_011110111001: DATA = 12'b100011011110;
            14'b11_011110111010: DATA = 12'b100011011011;
            14'b11_011110111011: DATA = 12'b100011011000;
            14'b11_011110111100: DATA = 12'b100011010101;
            14'b11_011110111101: DATA = 12'b100011010010;
            14'b11_011110111110: DATA = 12'b100011001110;
            14'b11_011110111111: DATA = 12'b100011001011;
            14'b11_011111000000: DATA = 12'b100011001000;
            14'b11_011111000001: DATA = 12'b100011000101;
            14'b11_011111000010: DATA = 12'b100011000010;
            14'b11_011111000011: DATA = 12'b100010111111;
            14'b11_011111000100: DATA = 12'b100010111100;
            14'b11_011111000101: DATA = 12'b100010111001;
            14'b11_011111000110: DATA = 12'b100010110101;
            14'b11_011111000111: DATA = 12'b100010110010;
            14'b11_011111001000: DATA = 12'b100010101111;
            14'b11_011111001001: DATA = 12'b100010101100;
            14'b11_011111001010: DATA = 12'b100010101001;
            14'b11_011111001011: DATA = 12'b100010100110;
            14'b11_011111001100: DATA = 12'b100010100011;
            14'b11_011111001101: DATA = 12'b100010011111;
            14'b11_011111001110: DATA = 12'b100010011100;
            14'b11_011111001111: DATA = 12'b100010011001;
            14'b11_011111010000: DATA = 12'b100010010110;
            14'b11_011111010001: DATA = 12'b100010010011;
            14'b11_011111010010: DATA = 12'b100010010000;
            14'b11_011111010011: DATA = 12'b100010001101;
            14'b11_011111010100: DATA = 12'b100010001010;
            14'b11_011111010101: DATA = 12'b100010000110;
            14'b11_011111010110: DATA = 12'b100010000011;
            14'b11_011111010111: DATA = 12'b100010000000;
            14'b11_011111011000: DATA = 12'b100001111101;
            14'b11_011111011001: DATA = 12'b100001111010;
            14'b11_011111011010: DATA = 12'b100001110111;
            14'b11_011111011011: DATA = 12'b100001110100;
            14'b11_011111011100: DATA = 12'b100001110000;
            14'b11_011111011101: DATA = 12'b100001101101;
            14'b11_011111011110: DATA = 12'b100001101010;
            14'b11_011111011111: DATA = 12'b100001100111;
            14'b11_011111100000: DATA = 12'b100001100100;
            14'b11_011111100001: DATA = 12'b100001100001;
            14'b11_011111100010: DATA = 12'b100001011110;
            14'b11_011111100011: DATA = 12'b100001011011;
            14'b11_011111100100: DATA = 12'b100001010111;
            14'b11_011111100101: DATA = 12'b100001010100;
            14'b11_011111100110: DATA = 12'b100001010001;
            14'b11_011111100111: DATA = 12'b100001001110;
            14'b11_011111101000: DATA = 12'b100001001011;
            14'b11_011111101001: DATA = 12'b100001001000;
            14'b11_011111101010: DATA = 12'b100001000101;
            14'b11_011111101011: DATA = 12'b100001000001;
            14'b11_011111101100: DATA = 12'b100000111110;
            14'b11_011111101101: DATA = 12'b100000111011;
            14'b11_011111101110: DATA = 12'b100000111000;
            14'b11_011111101111: DATA = 12'b100000110101;
            14'b11_011111110000: DATA = 12'b100000110010;
            14'b11_011111110001: DATA = 12'b100000101111;
            14'b11_011111110010: DATA = 12'b100000101011;
            14'b11_011111110011: DATA = 12'b100000101000;
            14'b11_011111110100: DATA = 12'b100000100101;
            14'b11_011111110101: DATA = 12'b100000100010;
            14'b11_011111110110: DATA = 12'b100000011111;
            14'b11_011111110111: DATA = 12'b100000011100;
            14'b11_011111111000: DATA = 12'b100000011001;
            14'b11_011111111001: DATA = 12'b100000010101;
            14'b11_011111111010: DATA = 12'b100000010010;
            14'b11_011111111011: DATA = 12'b100000001111;
            14'b11_011111111100: DATA = 12'b100000001100;
            14'b11_011111111101: DATA = 12'b100000001001;
            14'b11_011111111110: DATA = 12'b100000000110;
            14'b11_011111111111: DATA = 12'b100000000011;
            14'b11_100000000000: DATA = 12'b100000000000;
            14'b11_100000000001: DATA = 12'b100000000011;
            14'b11_100000000010: DATA = 12'b100000000110;
            14'b11_100000000011: DATA = 12'b100000001001;
            14'b11_100000000100: DATA = 12'b100000001100;
            14'b11_100000000101: DATA = 12'b100000001111;
            14'b11_100000000110: DATA = 12'b100000010010;
            14'b11_100000000111: DATA = 12'b100000010101;
            14'b11_100000001000: DATA = 12'b100000011001;
            14'b11_100000001001: DATA = 12'b100000011100;
            14'b11_100000001010: DATA = 12'b100000011111;
            14'b11_100000001011: DATA = 12'b100000100010;
            14'b11_100000001100: DATA = 12'b100000100101;
            14'b11_100000001101: DATA = 12'b100000101000;
            14'b11_100000001110: DATA = 12'b100000101011;
            14'b11_100000001111: DATA = 12'b100000101111;
            14'b11_100000010000: DATA = 12'b100000110010;
            14'b11_100000010001: DATA = 12'b100000110101;
            14'b11_100000010010: DATA = 12'b100000111000;
            14'b11_100000010011: DATA = 12'b100000111011;
            14'b11_100000010100: DATA = 12'b100000111110;
            14'b11_100000010101: DATA = 12'b100001000001;
            14'b11_100000010110: DATA = 12'b100001000101;
            14'b11_100000010111: DATA = 12'b100001001000;
            14'b11_100000011000: DATA = 12'b100001001011;
            14'b11_100000011001: DATA = 12'b100001001110;
            14'b11_100000011010: DATA = 12'b100001010001;
            14'b11_100000011011: DATA = 12'b100001010100;
            14'b11_100000011100: DATA = 12'b100001010111;
            14'b11_100000011101: DATA = 12'b100001011011;
            14'b11_100000011110: DATA = 12'b100001011110;
            14'b11_100000011111: DATA = 12'b100001100001;
            14'b11_100000100000: DATA = 12'b100001100100;
            14'b11_100000100001: DATA = 12'b100001100111;
            14'b11_100000100010: DATA = 12'b100001101010;
            14'b11_100000100011: DATA = 12'b100001101101;
            14'b11_100000100100: DATA = 12'b100001110000;
            14'b11_100000100101: DATA = 12'b100001110100;
            14'b11_100000100110: DATA = 12'b100001110111;
            14'b11_100000100111: DATA = 12'b100001111010;
            14'b11_100000101000: DATA = 12'b100001111101;
            14'b11_100000101001: DATA = 12'b100010000000;
            14'b11_100000101010: DATA = 12'b100010000011;
            14'b11_100000101011: DATA = 12'b100010000110;
            14'b11_100000101100: DATA = 12'b100010001010;
            14'b11_100000101101: DATA = 12'b100010001101;
            14'b11_100000101110: DATA = 12'b100010010000;
            14'b11_100000101111: DATA = 12'b100010010011;
            14'b11_100000110000: DATA = 12'b100010010110;
            14'b11_100000110001: DATA = 12'b100010011001;
            14'b11_100000110010: DATA = 12'b100010011100;
            14'b11_100000110011: DATA = 12'b100010011111;
            14'b11_100000110100: DATA = 12'b100010100011;
            14'b11_100000110101: DATA = 12'b100010100110;
            14'b11_100000110110: DATA = 12'b100010101001;
            14'b11_100000110111: DATA = 12'b100010101100;
            14'b11_100000111000: DATA = 12'b100010101111;
            14'b11_100000111001: DATA = 12'b100010110010;
            14'b11_100000111010: DATA = 12'b100010110101;
            14'b11_100000111011: DATA = 12'b100010111001;
            14'b11_100000111100: DATA = 12'b100010111100;
            14'b11_100000111101: DATA = 12'b100010111111;
            14'b11_100000111110: DATA = 12'b100011000010;
            14'b11_100000111111: DATA = 12'b100011000101;
            14'b11_100001000000: DATA = 12'b100011001000;
            14'b11_100001000001: DATA = 12'b100011001011;
            14'b11_100001000010: DATA = 12'b100011001110;
            14'b11_100001000011: DATA = 12'b100011010010;
            14'b11_100001000100: DATA = 12'b100011010101;
            14'b11_100001000101: DATA = 12'b100011011000;
            14'b11_100001000110: DATA = 12'b100011011011;
            14'b11_100001000111: DATA = 12'b100011011110;
            14'b11_100001001000: DATA = 12'b100011100001;
            14'b11_100001001001: DATA = 12'b100011100100;
            14'b11_100001001010: DATA = 12'b100011100111;
            14'b11_100001001011: DATA = 12'b100011101010;
            14'b11_100001001100: DATA = 12'b100011101110;
            14'b11_100001001101: DATA = 12'b100011110001;
            14'b11_100001001110: DATA = 12'b100011110100;
            14'b11_100001001111: DATA = 12'b100011110111;
            14'b11_100001010000: DATA = 12'b100011111010;
            14'b11_100001010001: DATA = 12'b100011111101;
            14'b11_100001010010: DATA = 12'b100100000000;
            14'b11_100001010011: DATA = 12'b100100000011;
            14'b11_100001010100: DATA = 12'b100100000111;
            14'b11_100001010101: DATA = 12'b100100001010;
            14'b11_100001010110: DATA = 12'b100100001101;
            14'b11_100001010111: DATA = 12'b100100010000;
            14'b11_100001011000: DATA = 12'b100100010011;
            14'b11_100001011001: DATA = 12'b100100010110;
            14'b11_100001011010: DATA = 12'b100100011001;
            14'b11_100001011011: DATA = 12'b100100011100;
            14'b11_100001011100: DATA = 12'b100100011111;
            14'b11_100001011101: DATA = 12'b100100100011;
            14'b11_100001011110: DATA = 12'b100100100110;
            14'b11_100001011111: DATA = 12'b100100101001;
            14'b11_100001100000: DATA = 12'b100100101100;
            14'b11_100001100001: DATA = 12'b100100101111;
            14'b11_100001100010: DATA = 12'b100100110010;
            14'b11_100001100011: DATA = 12'b100100110101;
            14'b11_100001100100: DATA = 12'b100100111000;
            14'b11_100001100101: DATA = 12'b100100111011;
            14'b11_100001100110: DATA = 12'b100100111110;
            14'b11_100001100111: DATA = 12'b100101000010;
            14'b11_100001101000: DATA = 12'b100101000101;
            14'b11_100001101001: DATA = 12'b100101001000;
            14'b11_100001101010: DATA = 12'b100101001011;
            14'b11_100001101011: DATA = 12'b100101001110;
            14'b11_100001101100: DATA = 12'b100101010001;
            14'b11_100001101101: DATA = 12'b100101010100;
            14'b11_100001101110: DATA = 12'b100101010111;
            14'b11_100001101111: DATA = 12'b100101011010;
            14'b11_100001110000: DATA = 12'b100101011101;
            14'b11_100001110001: DATA = 12'b100101100001;
            14'b11_100001110010: DATA = 12'b100101100100;
            14'b11_100001110011: DATA = 12'b100101100111;
            14'b11_100001110100: DATA = 12'b100101101010;
            14'b11_100001110101: DATA = 12'b100101101101;
            14'b11_100001110110: DATA = 12'b100101110000;
            14'b11_100001110111: DATA = 12'b100101110011;
            14'b11_100001111000: DATA = 12'b100101110110;
            14'b11_100001111001: DATA = 12'b100101111001;
            14'b11_100001111010: DATA = 12'b100101111100;
            14'b11_100001111011: DATA = 12'b100101111111;
            14'b11_100001111100: DATA = 12'b100110000011;
            14'b11_100001111101: DATA = 12'b100110000110;
            14'b11_100001111110: DATA = 12'b100110001001;
            14'b11_100001111111: DATA = 12'b100110001100;
            14'b11_100010000000: DATA = 12'b100110001111;
            14'b11_100010000001: DATA = 12'b100110010010;
            14'b11_100010000010: DATA = 12'b100110010101;
            14'b11_100010000011: DATA = 12'b100110011000;
            14'b11_100010000100: DATA = 12'b100110011011;
            14'b11_100010000101: DATA = 12'b100110011110;
            14'b11_100010000110: DATA = 12'b100110100001;
            14'b11_100010000111: DATA = 12'b100110100100;
            14'b11_100010001000: DATA = 12'b100110100111;
            14'b11_100010001001: DATA = 12'b100110101011;
            14'b11_100010001010: DATA = 12'b100110101110;
            14'b11_100010001011: DATA = 12'b100110110001;
            14'b11_100010001100: DATA = 12'b100110110100;
            14'b11_100010001101: DATA = 12'b100110110111;
            14'b11_100010001110: DATA = 12'b100110111010;
            14'b11_100010001111: DATA = 12'b100110111101;
            14'b11_100010010000: DATA = 12'b100111000000;
            14'b11_100010010001: DATA = 12'b100111000011;
            14'b11_100010010010: DATA = 12'b100111000110;
            14'b11_100010010011: DATA = 12'b100111001001;
            14'b11_100010010100: DATA = 12'b100111001100;
            14'b11_100010010101: DATA = 12'b100111001111;
            14'b11_100010010110: DATA = 12'b100111010010;
            14'b11_100010010111: DATA = 12'b100111010101;
            14'b11_100010011000: DATA = 12'b100111011000;
            14'b11_100010011001: DATA = 12'b100111011100;
            14'b11_100010011010: DATA = 12'b100111011111;
            14'b11_100010011011: DATA = 12'b100111100010;
            14'b11_100010011100: DATA = 12'b100111100101;
            14'b11_100010011101: DATA = 12'b100111101000;
            14'b11_100010011110: DATA = 12'b100111101011;
            14'b11_100010011111: DATA = 12'b100111101110;
            14'b11_100010100000: DATA = 12'b100111110001;
            14'b11_100010100001: DATA = 12'b100111110100;
            14'b11_100010100010: DATA = 12'b100111110111;
            14'b11_100010100011: DATA = 12'b100111111010;
            14'b11_100010100100: DATA = 12'b100111111101;
            14'b11_100010100101: DATA = 12'b101000000000;
            14'b11_100010100110: DATA = 12'b101000000011;
            14'b11_100010100111: DATA = 12'b101000000110;
            14'b11_100010101000: DATA = 12'b101000001001;
            14'b11_100010101001: DATA = 12'b101000001100;
            14'b11_100010101010: DATA = 12'b101000001111;
            14'b11_100010101011: DATA = 12'b101000010010;
            14'b11_100010101100: DATA = 12'b101000010101;
            14'b11_100010101101: DATA = 12'b101000011000;
            14'b11_100010101110: DATA = 12'b101000011011;
            14'b11_100010101111: DATA = 12'b101000011110;
            14'b11_100010110000: DATA = 12'b101000100001;
            14'b11_100010110001: DATA = 12'b101000100100;
            14'b11_100010110010: DATA = 12'b101000101000;
            14'b11_100010110011: DATA = 12'b101000101011;
            14'b11_100010110100: DATA = 12'b101000101110;
            14'b11_100010110101: DATA = 12'b101000110001;
            14'b11_100010110110: DATA = 12'b101000110100;
            14'b11_100010110111: DATA = 12'b101000110111;
            14'b11_100010111000: DATA = 12'b101000111010;
            14'b11_100010111001: DATA = 12'b101000111101;
            14'b11_100010111010: DATA = 12'b101001000000;
            14'b11_100010111011: DATA = 12'b101001000011;
            14'b11_100010111100: DATA = 12'b101001000110;
            14'b11_100010111101: DATA = 12'b101001001001;
            14'b11_100010111110: DATA = 12'b101001001100;
            14'b11_100010111111: DATA = 12'b101001001111;
            14'b11_100011000000: DATA = 12'b101001010010;
            14'b11_100011000001: DATA = 12'b101001010101;
            14'b11_100011000010: DATA = 12'b101001011000;
            14'b11_100011000011: DATA = 12'b101001011011;
            14'b11_100011000100: DATA = 12'b101001011110;
            14'b11_100011000101: DATA = 12'b101001100001;
            14'b11_100011000110: DATA = 12'b101001100100;
            14'b11_100011000111: DATA = 12'b101001100111;
            14'b11_100011001000: DATA = 12'b101001101010;
            14'b11_100011001001: DATA = 12'b101001101101;
            14'b11_100011001010: DATA = 12'b101001110000;
            14'b11_100011001011: DATA = 12'b101001110011;
            14'b11_100011001100: DATA = 12'b101001110110;
            14'b11_100011001101: DATA = 12'b101001111001;
            14'b11_100011001110: DATA = 12'b101001111100;
            14'b11_100011001111: DATA = 12'b101001111111;
            14'b11_100011010000: DATA = 12'b101010000010;
            14'b11_100011010001: DATA = 12'b101010000101;
            14'b11_100011010010: DATA = 12'b101010001000;
            14'b11_100011010011: DATA = 12'b101010001011;
            14'b11_100011010100: DATA = 12'b101010001110;
            14'b11_100011010101: DATA = 12'b101010010000;
            14'b11_100011010110: DATA = 12'b101010010011;
            14'b11_100011010111: DATA = 12'b101010010110;
            14'b11_100011011000: DATA = 12'b101010011001;
            14'b11_100011011001: DATA = 12'b101010011100;
            14'b11_100011011010: DATA = 12'b101010011111;
            14'b11_100011011011: DATA = 12'b101010100010;
            14'b11_100011011100: DATA = 12'b101010100101;
            14'b11_100011011101: DATA = 12'b101010101000;
            14'b11_100011011110: DATA = 12'b101010101011;
            14'b11_100011011111: DATA = 12'b101010101110;
            14'b11_100011100000: DATA = 12'b101010110001;
            14'b11_100011100001: DATA = 12'b101010110100;
            14'b11_100011100010: DATA = 12'b101010110111;
            14'b11_100011100011: DATA = 12'b101010111010;
            14'b11_100011100100: DATA = 12'b101010111101;
            14'b11_100011100101: DATA = 12'b101011000000;
            14'b11_100011100110: DATA = 12'b101011000011;
            14'b11_100011100111: DATA = 12'b101011000110;
            14'b11_100011101000: DATA = 12'b101011001001;
            14'b11_100011101001: DATA = 12'b101011001100;
            14'b11_100011101010: DATA = 12'b101011001111;
            14'b11_100011101011: DATA = 12'b101011010010;
            14'b11_100011101100: DATA = 12'b101011010100;
            14'b11_100011101101: DATA = 12'b101011010111;
            14'b11_100011101110: DATA = 12'b101011011010;
            14'b11_100011101111: DATA = 12'b101011011101;
            14'b11_100011110000: DATA = 12'b101011100000;
            14'b11_100011110001: DATA = 12'b101011100011;
            14'b11_100011110010: DATA = 12'b101011100110;
            14'b11_100011110011: DATA = 12'b101011101001;
            14'b11_100011110100: DATA = 12'b101011101100;
            14'b11_100011110101: DATA = 12'b101011101111;
            14'b11_100011110110: DATA = 12'b101011110010;
            14'b11_100011110111: DATA = 12'b101011110101;
            14'b11_100011111000: DATA = 12'b101011111000;
            14'b11_100011111001: DATA = 12'b101011111011;
            14'b11_100011111010: DATA = 12'b101011111101;
            14'b11_100011111011: DATA = 12'b101100000000;
            14'b11_100011111100: DATA = 12'b101100000011;
            14'b11_100011111101: DATA = 12'b101100000110;
            14'b11_100011111110: DATA = 12'b101100001001;
            14'b11_100011111111: DATA = 12'b101100001100;
            14'b11_100100000000: DATA = 12'b101100001111;
            14'b11_100100000001: DATA = 12'b101100010010;
            14'b11_100100000010: DATA = 12'b101100010101;
            14'b11_100100000011: DATA = 12'b101100011000;
            14'b11_100100000100: DATA = 12'b101100011010;
            14'b11_100100000101: DATA = 12'b101100011101;
            14'b11_100100000110: DATA = 12'b101100100000;
            14'b11_100100000111: DATA = 12'b101100100011;
            14'b11_100100001000: DATA = 12'b101100100110;
            14'b11_100100001001: DATA = 12'b101100101001;
            14'b11_100100001010: DATA = 12'b101100101100;
            14'b11_100100001011: DATA = 12'b101100101111;
            14'b11_100100001100: DATA = 12'b101100110010;
            14'b11_100100001101: DATA = 12'b101100110100;
            14'b11_100100001110: DATA = 12'b101100110111;
            14'b11_100100001111: DATA = 12'b101100111010;
            14'b11_100100010000: DATA = 12'b101100111101;
            14'b11_100100010001: DATA = 12'b101101000000;
            14'b11_100100010010: DATA = 12'b101101000011;
            14'b11_100100010011: DATA = 12'b101101000110;
            14'b11_100100010100: DATA = 12'b101101001000;
            14'b11_100100010101: DATA = 12'b101101001011;
            14'b11_100100010110: DATA = 12'b101101001110;
            14'b11_100100010111: DATA = 12'b101101010001;
            14'b11_100100011000: DATA = 12'b101101010100;
            14'b11_100100011001: DATA = 12'b101101010111;
            14'b11_100100011010: DATA = 12'b101101011010;
            14'b11_100100011011: DATA = 12'b101101011100;
            14'b11_100100011100: DATA = 12'b101101011111;
            14'b11_100100011101: DATA = 12'b101101100010;
            14'b11_100100011110: DATA = 12'b101101100101;
            14'b11_100100011111: DATA = 12'b101101101000;
            14'b11_100100100000: DATA = 12'b101101101011;
            14'b11_100100100001: DATA = 12'b101101101110;
            14'b11_100100100010: DATA = 12'b101101110000;
            14'b11_100100100011: DATA = 12'b101101110011;
            14'b11_100100100100: DATA = 12'b101101110110;
            14'b11_100100100101: DATA = 12'b101101111001;
            14'b11_100100100110: DATA = 12'b101101111100;
            14'b11_100100100111: DATA = 12'b101101111111;
            14'b11_100100101000: DATA = 12'b101110000001;
            14'b11_100100101001: DATA = 12'b101110000100;
            14'b11_100100101010: DATA = 12'b101110000111;
            14'b11_100100101011: DATA = 12'b101110001010;
            14'b11_100100101100: DATA = 12'b101110001101;
            14'b11_100100101101: DATA = 12'b101110001111;
            14'b11_100100101110: DATA = 12'b101110010010;
            14'b11_100100101111: DATA = 12'b101110010101;
            14'b11_100100110000: DATA = 12'b101110011000;
            14'b11_100100110001: DATA = 12'b101110011011;
            14'b11_100100110010: DATA = 12'b101110011101;
            14'b11_100100110011: DATA = 12'b101110100000;
            14'b11_100100110100: DATA = 12'b101110100011;
            14'b11_100100110101: DATA = 12'b101110100110;
            14'b11_100100110110: DATA = 12'b101110101001;
            14'b11_100100110111: DATA = 12'b101110101011;
            14'b11_100100111000: DATA = 12'b101110101110;
            14'b11_100100111001: DATA = 12'b101110110001;
            14'b11_100100111010: DATA = 12'b101110110100;
            14'b11_100100111011: DATA = 12'b101110110111;
            14'b11_100100111100: DATA = 12'b101110111001;
            14'b11_100100111101: DATA = 12'b101110111100;
            14'b11_100100111110: DATA = 12'b101110111111;
            14'b11_100100111111: DATA = 12'b101111000010;
            14'b11_100101000000: DATA = 12'b101111000100;
            14'b11_100101000001: DATA = 12'b101111000111;
            14'b11_100101000010: DATA = 12'b101111001010;
            14'b11_100101000011: DATA = 12'b101111001101;
            14'b11_100101000100: DATA = 12'b101111010000;
            14'b11_100101000101: DATA = 12'b101111010010;
            14'b11_100101000110: DATA = 12'b101111010101;
            14'b11_100101000111: DATA = 12'b101111011000;
            14'b11_100101001000: DATA = 12'b101111011011;
            14'b11_100101001001: DATA = 12'b101111011101;
            14'b11_100101001010: DATA = 12'b101111100000;
            14'b11_100101001011: DATA = 12'b101111100011;
            14'b11_100101001100: DATA = 12'b101111100110;
            14'b11_100101001101: DATA = 12'b101111101000;
            14'b11_100101001110: DATA = 12'b101111101011;
            14'b11_100101001111: DATA = 12'b101111101110;
            14'b11_100101010000: DATA = 12'b101111110000;
            14'b11_100101010001: DATA = 12'b101111110011;
            14'b11_100101010010: DATA = 12'b101111110110;
            14'b11_100101010011: DATA = 12'b101111111001;
            14'b11_100101010100: DATA = 12'b101111111011;
            14'b11_100101010101: DATA = 12'b101111111110;
            14'b11_100101010110: DATA = 12'b110000000001;
            14'b11_100101010111: DATA = 12'b110000000100;
            14'b11_100101011000: DATA = 12'b110000000110;
            14'b11_100101011001: DATA = 12'b110000001001;
            14'b11_100101011010: DATA = 12'b110000001100;
            14'b11_100101011011: DATA = 12'b110000001110;
            14'b11_100101011100: DATA = 12'b110000010001;
            14'b11_100101011101: DATA = 12'b110000010100;
            14'b11_100101011110: DATA = 12'b110000010110;
            14'b11_100101011111: DATA = 12'b110000011001;
            14'b11_100101100000: DATA = 12'b110000011100;
            14'b11_100101100001: DATA = 12'b110000011111;
            14'b11_100101100010: DATA = 12'b110000100001;
            14'b11_100101100011: DATA = 12'b110000100100;
            14'b11_100101100100: DATA = 12'b110000100111;
            14'b11_100101100101: DATA = 12'b110000101001;
            14'b11_100101100110: DATA = 12'b110000101100;
            14'b11_100101100111: DATA = 12'b110000101111;
            14'b11_100101101000: DATA = 12'b110000110001;
            14'b11_100101101001: DATA = 12'b110000110100;
            14'b11_100101101010: DATA = 12'b110000110111;
            14'b11_100101101011: DATA = 12'b110000111001;
            14'b11_100101101100: DATA = 12'b110000111100;
            14'b11_100101101101: DATA = 12'b110000111111;
            14'b11_100101101110: DATA = 12'b110001000001;
            14'b11_100101101111: DATA = 12'b110001000100;
            14'b11_100101110000: DATA = 12'b110001000111;
            14'b11_100101110001: DATA = 12'b110001001001;
            14'b11_100101110010: DATA = 12'b110001001100;
            14'b11_100101110011: DATA = 12'b110001001111;
            14'b11_100101110100: DATA = 12'b110001010001;
            14'b11_100101110101: DATA = 12'b110001010100;
            14'b11_100101110110: DATA = 12'b110001010111;
            14'b11_100101110111: DATA = 12'b110001011001;
            14'b11_100101111000: DATA = 12'b110001011100;
            14'b11_100101111001: DATA = 12'b110001011110;
            14'b11_100101111010: DATA = 12'b110001100001;
            14'b11_100101111011: DATA = 12'b110001100100;
            14'b11_100101111100: DATA = 12'b110001100110;
            14'b11_100101111101: DATA = 12'b110001101001;
            14'b11_100101111110: DATA = 12'b110001101100;
            14'b11_100101111111: DATA = 12'b110001101110;
            14'b11_100110000000: DATA = 12'b110001110001;
            14'b11_100110000001: DATA = 12'b110001110011;
            14'b11_100110000010: DATA = 12'b110001110110;
            14'b11_100110000011: DATA = 12'b110001111001;
            14'b11_100110000100: DATA = 12'b110001111011;
            14'b11_100110000101: DATA = 12'b110001111110;
            14'b11_100110000110: DATA = 12'b110010000000;
            14'b11_100110000111: DATA = 12'b110010000011;
            14'b11_100110001000: DATA = 12'b110010000110;
            14'b11_100110001001: DATA = 12'b110010001000;
            14'b11_100110001010: DATA = 12'b110010001011;
            14'b11_100110001011: DATA = 12'b110010001101;
            14'b11_100110001100: DATA = 12'b110010010000;
            14'b11_100110001101: DATA = 12'b110010010010;
            14'b11_100110001110: DATA = 12'b110010010101;
            14'b11_100110001111: DATA = 12'b110010011000;
            14'b11_100110010000: DATA = 12'b110010011010;
            14'b11_100110010001: DATA = 12'b110010011101;
            14'b11_100110010010: DATA = 12'b110010011111;
            14'b11_100110010011: DATA = 12'b110010100010;
            14'b11_100110010100: DATA = 12'b110010100100;
            14'b11_100110010101: DATA = 12'b110010100111;
            14'b11_100110010110: DATA = 12'b110010101010;
            14'b11_100110010111: DATA = 12'b110010101100;
            14'b11_100110011000: DATA = 12'b110010101111;
            14'b11_100110011001: DATA = 12'b110010110001;
            14'b11_100110011010: DATA = 12'b110010110100;
            14'b11_100110011011: DATA = 12'b110010110110;
            14'b11_100110011100: DATA = 12'b110010111001;
            14'b11_100110011101: DATA = 12'b110010111011;
            14'b11_100110011110: DATA = 12'b110010111110;
            14'b11_100110011111: DATA = 12'b110011000000;
            14'b11_100110100000: DATA = 12'b110011000011;
            14'b11_100110100001: DATA = 12'b110011000101;
            14'b11_100110100010: DATA = 12'b110011001000;
            14'b11_100110100011: DATA = 12'b110011001010;
            14'b11_100110100100: DATA = 12'b110011001101;
            14'b11_100110100101: DATA = 12'b110011001111;
            14'b11_100110100110: DATA = 12'b110011010010;
            14'b11_100110100111: DATA = 12'b110011010100;
            14'b11_100110101000: DATA = 12'b110011010111;
            14'b11_100110101001: DATA = 12'b110011011001;
            14'b11_100110101010: DATA = 12'b110011011100;
            14'b11_100110101011: DATA = 12'b110011011110;
            14'b11_100110101100: DATA = 12'b110011100001;
            14'b11_100110101101: DATA = 12'b110011100011;
            14'b11_100110101110: DATA = 12'b110011100110;
            14'b11_100110101111: DATA = 12'b110011101000;
            14'b11_100110110000: DATA = 12'b110011101011;
            14'b11_100110110001: DATA = 12'b110011101101;
            14'b11_100110110010: DATA = 12'b110011110000;
            14'b11_100110110011: DATA = 12'b110011110010;
            14'b11_100110110100: DATA = 12'b110011110101;
            14'b11_100110110101: DATA = 12'b110011110111;
            14'b11_100110110110: DATA = 12'b110011111010;
            14'b11_100110110111: DATA = 12'b110011111100;
            14'b11_100110111000: DATA = 12'b110011111111;
            14'b11_100110111001: DATA = 12'b110100000001;
            14'b11_100110111010: DATA = 12'b110100000011;
            14'b11_100110111011: DATA = 12'b110100000110;
            14'b11_100110111100: DATA = 12'b110100001000;
            14'b11_100110111101: DATA = 12'b110100001011;
            14'b11_100110111110: DATA = 12'b110100001101;
            14'b11_100110111111: DATA = 12'b110100010000;
            14'b11_100111000000: DATA = 12'b110100010010;
            14'b11_100111000001: DATA = 12'b110100010101;
            14'b11_100111000010: DATA = 12'b110100010111;
            14'b11_100111000011: DATA = 12'b110100011001;
            14'b11_100111000100: DATA = 12'b110100011100;
            14'b11_100111000101: DATA = 12'b110100011110;
            14'b11_100111000110: DATA = 12'b110100100001;
            14'b11_100111000111: DATA = 12'b110100100011;
            14'b11_100111001000: DATA = 12'b110100100101;
            14'b11_100111001001: DATA = 12'b110100101000;
            14'b11_100111001010: DATA = 12'b110100101010;
            14'b11_100111001011: DATA = 12'b110100101101;
            14'b11_100111001100: DATA = 12'b110100101111;
            14'b11_100111001101: DATA = 12'b110100110001;
            14'b11_100111001110: DATA = 12'b110100110100;
            14'b11_100111001111: DATA = 12'b110100110110;
            14'b11_100111010000: DATA = 12'b110100111001;
            14'b11_100111010001: DATA = 12'b110100111011;
            14'b11_100111010010: DATA = 12'b110100111101;
            14'b11_100111010011: DATA = 12'b110101000000;
            14'b11_100111010100: DATA = 12'b110101000010;
            14'b11_100111010101: DATA = 12'b110101000100;
            14'b11_100111010110: DATA = 12'b110101000111;
            14'b11_100111010111: DATA = 12'b110101001001;
            14'b11_100111011000: DATA = 12'b110101001011;
            14'b11_100111011001: DATA = 12'b110101001110;
            14'b11_100111011010: DATA = 12'b110101010000;
            14'b11_100111011011: DATA = 12'b110101010011;
            14'b11_100111011100: DATA = 12'b110101010101;
            14'b11_100111011101: DATA = 12'b110101010111;
            14'b11_100111011110: DATA = 12'b110101011010;
            14'b11_100111011111: DATA = 12'b110101011100;
            14'b11_100111100000: DATA = 12'b110101011110;
            14'b11_100111100001: DATA = 12'b110101100001;
            14'b11_100111100010: DATA = 12'b110101100011;
            14'b11_100111100011: DATA = 12'b110101100101;
            14'b11_100111100100: DATA = 12'b110101100111;
            14'b11_100111100101: DATA = 12'b110101101010;
            14'b11_100111100110: DATA = 12'b110101101100;
            14'b11_100111100111: DATA = 12'b110101101110;
            14'b11_100111101000: DATA = 12'b110101110001;
            14'b11_100111101001: DATA = 12'b110101110011;
            14'b11_100111101010: DATA = 12'b110101110101;
            14'b11_100111101011: DATA = 12'b110101111000;
            14'b11_100111101100: DATA = 12'b110101111010;
            14'b11_100111101101: DATA = 12'b110101111100;
            14'b11_100111101110: DATA = 12'b110101111110;
            14'b11_100111101111: DATA = 12'b110110000001;
            14'b11_100111110000: DATA = 12'b110110000011;
            14'b11_100111110001: DATA = 12'b110110000101;
            14'b11_100111110010: DATA = 12'b110110001000;
            14'b11_100111110011: DATA = 12'b110110001010;
            14'b11_100111110100: DATA = 12'b110110001100;
            14'b11_100111110101: DATA = 12'b110110001110;
            14'b11_100111110110: DATA = 12'b110110010001;
            14'b11_100111110111: DATA = 12'b110110010011;
            14'b11_100111111000: DATA = 12'b110110010101;
            14'b11_100111111001: DATA = 12'b110110010111;
            14'b11_100111111010: DATA = 12'b110110011010;
            14'b11_100111111011: DATA = 12'b110110011100;
            14'b11_100111111100: DATA = 12'b110110011110;
            14'b11_100111111101: DATA = 12'b110110100000;
            14'b11_100111111110: DATA = 12'b110110100011;
            14'b11_100111111111: DATA = 12'b110110100101;
            14'b11_101000000000: DATA = 12'b110110100111;
            14'b11_101000000001: DATA = 12'b110110101001;
            14'b11_101000000010: DATA = 12'b110110101011;
            14'b11_101000000011: DATA = 12'b110110101110;
            14'b11_101000000100: DATA = 12'b110110110000;
            14'b11_101000000101: DATA = 12'b110110110010;
            14'b11_101000000110: DATA = 12'b110110110100;
            14'b11_101000000111: DATA = 12'b110110110110;
            14'b11_101000001000: DATA = 12'b110110111001;
            14'b11_101000001001: DATA = 12'b110110111011;
            14'b11_101000001010: DATA = 12'b110110111101;
            14'b11_101000001011: DATA = 12'b110110111111;
            14'b11_101000001100: DATA = 12'b110111000001;
            14'b11_101000001101: DATA = 12'b110111000100;
            14'b11_101000001110: DATA = 12'b110111000110;
            14'b11_101000001111: DATA = 12'b110111001000;
            14'b11_101000010000: DATA = 12'b110111001010;
            14'b11_101000010001: DATA = 12'b110111001100;
            14'b11_101000010010: DATA = 12'b110111001110;
            14'b11_101000010011: DATA = 12'b110111010001;
            14'b11_101000010100: DATA = 12'b110111010011;
            14'b11_101000010101: DATA = 12'b110111010101;
            14'b11_101000010110: DATA = 12'b110111010111;
            14'b11_101000010111: DATA = 12'b110111011001;
            14'b11_101000011000: DATA = 12'b110111011011;
            14'b11_101000011001: DATA = 12'b110111011101;
            14'b11_101000011010: DATA = 12'b110111100000;
            14'b11_101000011011: DATA = 12'b110111100010;
            14'b11_101000011100: DATA = 12'b110111100100;
            14'b11_101000011101: DATA = 12'b110111100110;
            14'b11_101000011110: DATA = 12'b110111101000;
            14'b11_101000011111: DATA = 12'b110111101010;
            14'b11_101000100000: DATA = 12'b110111101100;
            14'b11_101000100001: DATA = 12'b110111101110;
            14'b11_101000100010: DATA = 12'b110111110000;
            14'b11_101000100011: DATA = 12'b110111110011;
            14'b11_101000100100: DATA = 12'b110111110101;
            14'b11_101000100101: DATA = 12'b110111110111;
            14'b11_101000100110: DATA = 12'b110111111001;
            14'b11_101000100111: DATA = 12'b110111111011;
            14'b11_101000101000: DATA = 12'b110111111101;
            14'b11_101000101001: DATA = 12'b110111111111;
            14'b11_101000101010: DATA = 12'b111000000001;
            14'b11_101000101011: DATA = 12'b111000000011;
            14'b11_101000101100: DATA = 12'b111000000101;
            14'b11_101000101101: DATA = 12'b111000000111;
            14'b11_101000101110: DATA = 12'b111000001001;
            14'b11_101000101111: DATA = 12'b111000001011;
            14'b11_101000110000: DATA = 12'b111000001110;
            14'b11_101000110001: DATA = 12'b111000010000;
            14'b11_101000110010: DATA = 12'b111000010010;
            14'b11_101000110011: DATA = 12'b111000010100;
            14'b11_101000110100: DATA = 12'b111000010110;
            14'b11_101000110101: DATA = 12'b111000011000;
            14'b11_101000110110: DATA = 12'b111000011010;
            14'b11_101000110111: DATA = 12'b111000011100;
            14'b11_101000111000: DATA = 12'b111000011110;
            14'b11_101000111001: DATA = 12'b111000100000;
            14'b11_101000111010: DATA = 12'b111000100010;
            14'b11_101000111011: DATA = 12'b111000100100;
            14'b11_101000111100: DATA = 12'b111000100110;
            14'b11_101000111101: DATA = 12'b111000101000;
            14'b11_101000111110: DATA = 12'b111000101010;
            14'b11_101000111111: DATA = 12'b111000101100;
            14'b11_101001000000: DATA = 12'b111000101110;
            14'b11_101001000001: DATA = 12'b111000110000;
            14'b11_101001000010: DATA = 12'b111000110010;
            14'b11_101001000011: DATA = 12'b111000110100;
            14'b11_101001000100: DATA = 12'b111000110110;
            14'b11_101001000101: DATA = 12'b111000111000;
            14'b11_101001000110: DATA = 12'b111000111010;
            14'b11_101001000111: DATA = 12'b111000111100;
            14'b11_101001001000: DATA = 12'b111000111110;
            14'b11_101001001001: DATA = 12'b111001000000;
            14'b11_101001001010: DATA = 12'b111001000010;
            14'b11_101001001011: DATA = 12'b111001000100;
            14'b11_101001001100: DATA = 12'b111001000101;
            14'b11_101001001101: DATA = 12'b111001000111;
            14'b11_101001001110: DATA = 12'b111001001001;
            14'b11_101001001111: DATA = 12'b111001001011;
            14'b11_101001010000: DATA = 12'b111001001101;
            14'b11_101001010001: DATA = 12'b111001001111;
            14'b11_101001010010: DATA = 12'b111001010001;
            14'b11_101001010011: DATA = 12'b111001010011;
            14'b11_101001010100: DATA = 12'b111001010101;
            14'b11_101001010101: DATA = 12'b111001010111;
            14'b11_101001010110: DATA = 12'b111001011001;
            14'b11_101001010111: DATA = 12'b111001011011;
            14'b11_101001011000: DATA = 12'b111001011101;
            14'b11_101001011001: DATA = 12'b111001011110;
            14'b11_101001011010: DATA = 12'b111001100000;
            14'b11_101001011011: DATA = 12'b111001100010;
            14'b11_101001011100: DATA = 12'b111001100100;
            14'b11_101001011101: DATA = 12'b111001100110;
            14'b11_101001011110: DATA = 12'b111001101000;
            14'b11_101001011111: DATA = 12'b111001101010;
            14'b11_101001100000: DATA = 12'b111001101100;
            14'b11_101001100001: DATA = 12'b111001101110;
            14'b11_101001100010: DATA = 12'b111001101111;
            14'b11_101001100011: DATA = 12'b111001110001;
            14'b11_101001100100: DATA = 12'b111001110011;
            14'b11_101001100101: DATA = 12'b111001110101;
            14'b11_101001100110: DATA = 12'b111001110111;
            14'b11_101001100111: DATA = 12'b111001111001;
            14'b11_101001101000: DATA = 12'b111001111011;
            14'b11_101001101001: DATA = 12'b111001111100;
            14'b11_101001101010: DATA = 12'b111001111110;
            14'b11_101001101011: DATA = 12'b111010000000;
            14'b11_101001101100: DATA = 12'b111010000010;
            14'b11_101001101101: DATA = 12'b111010000100;
            14'b11_101001101110: DATA = 12'b111010000101;
            14'b11_101001101111: DATA = 12'b111010000111;
            14'b11_101001110000: DATA = 12'b111010001001;
            14'b11_101001110001: DATA = 12'b111010001011;
            14'b11_101001110010: DATA = 12'b111010001101;
            14'b11_101001110011: DATA = 12'b111010001111;
            14'b11_101001110100: DATA = 12'b111010010000;
            14'b11_101001110101: DATA = 12'b111010010010;
            14'b11_101001110110: DATA = 12'b111010010100;
            14'b11_101001110111: DATA = 12'b111010010110;
            14'b11_101001111000: DATA = 12'b111010010111;
            14'b11_101001111001: DATA = 12'b111010011001;
            14'b11_101001111010: DATA = 12'b111010011011;
            14'b11_101001111011: DATA = 12'b111010011101;
            14'b11_101001111100: DATA = 12'b111010011111;
            14'b11_101001111101: DATA = 12'b111010100000;
            14'b11_101001111110: DATA = 12'b111010100010;
            14'b11_101001111111: DATA = 12'b111010100100;
            14'b11_101010000000: DATA = 12'b111010100110;
            14'b11_101010000001: DATA = 12'b111010100111;
            14'b11_101010000010: DATA = 12'b111010101001;
            14'b11_101010000011: DATA = 12'b111010101011;
            14'b11_101010000100: DATA = 12'b111010101100;
            14'b11_101010000101: DATA = 12'b111010101110;
            14'b11_101010000110: DATA = 12'b111010110000;
            14'b11_101010000111: DATA = 12'b111010110010;
            14'b11_101010001000: DATA = 12'b111010110011;
            14'b11_101010001001: DATA = 12'b111010110101;
            14'b11_101010001010: DATA = 12'b111010110111;
            14'b11_101010001011: DATA = 12'b111010111000;
            14'b11_101010001100: DATA = 12'b111010111010;
            14'b11_101010001101: DATA = 12'b111010111100;
            14'b11_101010001110: DATA = 12'b111010111110;
            14'b11_101010001111: DATA = 12'b111010111111;
            14'b11_101010010000: DATA = 12'b111011000001;
            14'b11_101010010001: DATA = 12'b111011000011;
            14'b11_101010010010: DATA = 12'b111011000100;
            14'b11_101010010011: DATA = 12'b111011000110;
            14'b11_101010010100: DATA = 12'b111011001000;
            14'b11_101010010101: DATA = 12'b111011001001;
            14'b11_101010010110: DATA = 12'b111011001011;
            14'b11_101010010111: DATA = 12'b111011001101;
            14'b11_101010011000: DATA = 12'b111011001110;
            14'b11_101010011001: DATA = 12'b111011010000;
            14'b11_101010011010: DATA = 12'b111011010010;
            14'b11_101010011011: DATA = 12'b111011010011;
            14'b11_101010011100: DATA = 12'b111011010101;
            14'b11_101010011101: DATA = 12'b111011010110;
            14'b11_101010011110: DATA = 12'b111011011000;
            14'b11_101010011111: DATA = 12'b111011011010;
            14'b11_101010100000: DATA = 12'b111011011011;
            14'b11_101010100001: DATA = 12'b111011011101;
            14'b11_101010100010: DATA = 12'b111011011110;
            14'b11_101010100011: DATA = 12'b111011100000;
            14'b11_101010100100: DATA = 12'b111011100010;
            14'b11_101010100101: DATA = 12'b111011100011;
            14'b11_101010100110: DATA = 12'b111011100101;
            14'b11_101010100111: DATA = 12'b111011100110;
            14'b11_101010101000: DATA = 12'b111011101000;
            14'b11_101010101001: DATA = 12'b111011101010;
            14'b11_101010101010: DATA = 12'b111011101011;
            14'b11_101010101011: DATA = 12'b111011101101;
            14'b11_101010101100: DATA = 12'b111011101110;
            14'b11_101010101101: DATA = 12'b111011110000;
            14'b11_101010101110: DATA = 12'b111011110001;
            14'b11_101010101111: DATA = 12'b111011110011;
            14'b11_101010110000: DATA = 12'b111011110101;
            14'b11_101010110001: DATA = 12'b111011110110;
            14'b11_101010110010: DATA = 12'b111011111000;
            14'b11_101010110011: DATA = 12'b111011111001;
            14'b11_101010110100: DATA = 12'b111011111011;
            14'b11_101010110101: DATA = 12'b111011111100;
            14'b11_101010110110: DATA = 12'b111011111110;
            14'b11_101010110111: DATA = 12'b111011111111;
            14'b11_101010111000: DATA = 12'b111100000001;
            14'b11_101010111001: DATA = 12'b111100000010;
            14'b11_101010111010: DATA = 12'b111100000100;
            14'b11_101010111011: DATA = 12'b111100000101;
            14'b11_101010111100: DATA = 12'b111100000111;
            14'b11_101010111101: DATA = 12'b111100001000;
            14'b11_101010111110: DATA = 12'b111100001010;
            14'b11_101010111111: DATA = 12'b111100001011;
            14'b11_101011000000: DATA = 12'b111100001101;
            14'b11_101011000001: DATA = 12'b111100001110;
            14'b11_101011000010: DATA = 12'b111100010000;
            14'b11_101011000011: DATA = 12'b111100010001;
            14'b11_101011000100: DATA = 12'b111100010011;
            14'b11_101011000101: DATA = 12'b111100010100;
            14'b11_101011000110: DATA = 12'b111100010110;
            14'b11_101011000111: DATA = 12'b111100010111;
            14'b11_101011001000: DATA = 12'b111100011000;
            14'b11_101011001001: DATA = 12'b111100011010;
            14'b11_101011001010: DATA = 12'b111100011011;
            14'b11_101011001011: DATA = 12'b111100011101;
            14'b11_101011001100: DATA = 12'b111100011110;
            14'b11_101011001101: DATA = 12'b111100100000;
            14'b11_101011001110: DATA = 12'b111100100001;
            14'b11_101011001111: DATA = 12'b111100100011;
            14'b11_101011010000: DATA = 12'b111100100100;
            14'b11_101011010001: DATA = 12'b111100100101;
            14'b11_101011010010: DATA = 12'b111100100111;
            14'b11_101011010011: DATA = 12'b111100101000;
            14'b11_101011010100: DATA = 12'b111100101010;
            14'b11_101011010101: DATA = 12'b111100101011;
            14'b11_101011010110: DATA = 12'b111100101100;
            14'b11_101011010111: DATA = 12'b111100101110;
            14'b11_101011011000: DATA = 12'b111100101111;
            14'b11_101011011001: DATA = 12'b111100110000;
            14'b11_101011011010: DATA = 12'b111100110010;
            14'b11_101011011011: DATA = 12'b111100110011;
            14'b11_101011011100: DATA = 12'b111100110101;
            14'b11_101011011101: DATA = 12'b111100110110;
            14'b11_101011011110: DATA = 12'b111100110111;
            14'b11_101011011111: DATA = 12'b111100111001;
            14'b11_101011100000: DATA = 12'b111100111010;
            14'b11_101011100001: DATA = 12'b111100111011;
            14'b11_101011100010: DATA = 12'b111100111101;
            14'b11_101011100011: DATA = 12'b111100111110;
            14'b11_101011100100: DATA = 12'b111100111111;
            14'b11_101011100101: DATA = 12'b111101000001;
            14'b11_101011100110: DATA = 12'b111101000010;
            14'b11_101011100111: DATA = 12'b111101000011;
            14'b11_101011101000: DATA = 12'b111101000101;
            14'b11_101011101001: DATA = 12'b111101000110;
            14'b11_101011101010: DATA = 12'b111101000111;
            14'b11_101011101011: DATA = 12'b111101001000;
            14'b11_101011101100: DATA = 12'b111101001010;
            14'b11_101011101101: DATA = 12'b111101001011;
            14'b11_101011101110: DATA = 12'b111101001100;
            14'b11_101011101111: DATA = 12'b111101001110;
            14'b11_101011110000: DATA = 12'b111101001111;
            14'b11_101011110001: DATA = 12'b111101010000;
            14'b11_101011110010: DATA = 12'b111101010001;
            14'b11_101011110011: DATA = 12'b111101010011;
            14'b11_101011110100: DATA = 12'b111101010100;
            14'b11_101011110101: DATA = 12'b111101010101;
            14'b11_101011110110: DATA = 12'b111101010110;
            14'b11_101011110111: DATA = 12'b111101011000;
            14'b11_101011111000: DATA = 12'b111101011001;
            14'b11_101011111001: DATA = 12'b111101011010;
            14'b11_101011111010: DATA = 12'b111101011011;
            14'b11_101011111011: DATA = 12'b111101011101;
            14'b11_101011111100: DATA = 12'b111101011110;
            14'b11_101011111101: DATA = 12'b111101011111;
            14'b11_101011111110: DATA = 12'b111101100000;
            14'b11_101011111111: DATA = 12'b111101100001;
            14'b11_101100000000: DATA = 12'b111101100011;
            14'b11_101100000001: DATA = 12'b111101100100;
            14'b11_101100000010: DATA = 12'b111101100101;
            14'b11_101100000011: DATA = 12'b111101100110;
            14'b11_101100000100: DATA = 12'b111101100111;
            14'b11_101100000101: DATA = 12'b111101101001;
            14'b11_101100000110: DATA = 12'b111101101010;
            14'b11_101100000111: DATA = 12'b111101101011;
            14'b11_101100001000: DATA = 12'b111101101100;
            14'b11_101100001001: DATA = 12'b111101101101;
            14'b11_101100001010: DATA = 12'b111101101110;
            14'b11_101100001011: DATA = 12'b111101110000;
            14'b11_101100001100: DATA = 12'b111101110001;
            14'b11_101100001101: DATA = 12'b111101110010;
            14'b11_101100001110: DATA = 12'b111101110011;
            14'b11_101100001111: DATA = 12'b111101110100;
            14'b11_101100010000: DATA = 12'b111101110101;
            14'b11_101100010001: DATA = 12'b111101110110;
            14'b11_101100010010: DATA = 12'b111101111000;
            14'b11_101100010011: DATA = 12'b111101111001;
            14'b11_101100010100: DATA = 12'b111101111010;
            14'b11_101100010101: DATA = 12'b111101111011;
            14'b11_101100010110: DATA = 12'b111101111100;
            14'b11_101100010111: DATA = 12'b111101111101;
            14'b11_101100011000: DATA = 12'b111101111110;
            14'b11_101100011001: DATA = 12'b111101111111;
            14'b11_101100011010: DATA = 12'b111110000000;
            14'b11_101100011011: DATA = 12'b111110000001;
            14'b11_101100011100: DATA = 12'b111110000011;
            14'b11_101100011101: DATA = 12'b111110000100;
            14'b11_101100011110: DATA = 12'b111110000101;
            14'b11_101100011111: DATA = 12'b111110000110;
            14'b11_101100100000: DATA = 12'b111110000111;
            14'b11_101100100001: DATA = 12'b111110001000;
            14'b11_101100100010: DATA = 12'b111110001001;
            14'b11_101100100011: DATA = 12'b111110001010;
            14'b11_101100100100: DATA = 12'b111110001011;
            14'b11_101100100101: DATA = 12'b111110001100;
            14'b11_101100100110: DATA = 12'b111110001101;
            14'b11_101100100111: DATA = 12'b111110001110;
            14'b11_101100101000: DATA = 12'b111110001111;
            14'b11_101100101001: DATA = 12'b111110010000;
            14'b11_101100101010: DATA = 12'b111110010001;
            14'b11_101100101011: DATA = 12'b111110010010;
            14'b11_101100101100: DATA = 12'b111110010011;
            14'b11_101100101101: DATA = 12'b111110010100;
            14'b11_101100101110: DATA = 12'b111110010101;
            14'b11_101100101111: DATA = 12'b111110010110;
            14'b11_101100110000: DATA = 12'b111110010111;
            14'b11_101100110001: DATA = 12'b111110011000;
            14'b11_101100110010: DATA = 12'b111110011001;
            14'b11_101100110011: DATA = 12'b111110011010;
            14'b11_101100110100: DATA = 12'b111110011011;
            14'b11_101100110101: DATA = 12'b111110011100;
            14'b11_101100110110: DATA = 12'b111110011101;
            14'b11_101100110111: DATA = 12'b111110011110;
            14'b11_101100111000: DATA = 12'b111110011111;
            14'b11_101100111001: DATA = 12'b111110100000;
            14'b11_101100111010: DATA = 12'b111110100001;
            14'b11_101100111011: DATA = 12'b111110100010;
            14'b11_101100111100: DATA = 12'b111110100011;
            14'b11_101100111101: DATA = 12'b111110100100;
            14'b11_101100111110: DATA = 12'b111110100101;
            14'b11_101100111111: DATA = 12'b111110100101;
            14'b11_101101000000: DATA = 12'b111110100110;
            14'b11_101101000001: DATA = 12'b111110100111;
            14'b11_101101000010: DATA = 12'b111110101000;
            14'b11_101101000011: DATA = 12'b111110101001;
            14'b11_101101000100: DATA = 12'b111110101010;
            14'b11_101101000101: DATA = 12'b111110101011;
            14'b11_101101000110: DATA = 12'b111110101100;
            14'b11_101101000111: DATA = 12'b111110101101;
            14'b11_101101001000: DATA = 12'b111110101110;
            14'b11_101101001001: DATA = 12'b111110101110;
            14'b11_101101001010: DATA = 12'b111110101111;
            14'b11_101101001011: DATA = 12'b111110110000;
            14'b11_101101001100: DATA = 12'b111110110001;
            14'b11_101101001101: DATA = 12'b111110110010;
            14'b11_101101001110: DATA = 12'b111110110011;
            14'b11_101101001111: DATA = 12'b111110110100;
            14'b11_101101010000: DATA = 12'b111110110100;
            14'b11_101101010001: DATA = 12'b111110110101;
            14'b11_101101010010: DATA = 12'b111110110110;
            14'b11_101101010011: DATA = 12'b111110110111;
            14'b11_101101010100: DATA = 12'b111110111000;
            14'b11_101101010101: DATA = 12'b111110111000;
            14'b11_101101010110: DATA = 12'b111110111001;
            14'b11_101101010111: DATA = 12'b111110111010;
            14'b11_101101011000: DATA = 12'b111110111011;
            14'b11_101101011001: DATA = 12'b111110111100;
            14'b11_101101011010: DATA = 12'b111110111100;
            14'b11_101101011011: DATA = 12'b111110111101;
            14'b11_101101011100: DATA = 12'b111110111110;
            14'b11_101101011101: DATA = 12'b111110111111;
            14'b11_101101011110: DATA = 12'b111111000000;
            14'b11_101101011111: DATA = 12'b111111000000;
            14'b11_101101100000: DATA = 12'b111111000001;
            14'b11_101101100001: DATA = 12'b111111000010;
            14'b11_101101100010: DATA = 12'b111111000011;
            14'b11_101101100011: DATA = 12'b111111000011;
            14'b11_101101100100: DATA = 12'b111111000100;
            14'b11_101101100101: DATA = 12'b111111000101;
            14'b11_101101100110: DATA = 12'b111111000110;
            14'b11_101101100111: DATA = 12'b111111000110;
            14'b11_101101101000: DATA = 12'b111111000111;
            14'b11_101101101001: DATA = 12'b111111001000;
            14'b11_101101101010: DATA = 12'b111111001001;
            14'b11_101101101011: DATA = 12'b111111001001;
            14'b11_101101101100: DATA = 12'b111111001010;
            14'b11_101101101101: DATA = 12'b111111001011;
            14'b11_101101101110: DATA = 12'b111111001011;
            14'b11_101101101111: DATA = 12'b111111001100;
            14'b11_101101110000: DATA = 12'b111111001101;
            14'b11_101101110001: DATA = 12'b111111001101;
            14'b11_101101110010: DATA = 12'b111111001110;
            14'b11_101101110011: DATA = 12'b111111001111;
            14'b11_101101110100: DATA = 12'b111111001111;
            14'b11_101101110101: DATA = 12'b111111010000;
            14'b11_101101110110: DATA = 12'b111111010001;
            14'b11_101101110111: DATA = 12'b111111010001;
            14'b11_101101111000: DATA = 12'b111111010010;
            14'b11_101101111001: DATA = 12'b111111010011;
            14'b11_101101111010: DATA = 12'b111111010011;
            14'b11_101101111011: DATA = 12'b111111010100;
            14'b11_101101111100: DATA = 12'b111111010101;
            14'b11_101101111101: DATA = 12'b111111010101;
            14'b11_101101111110: DATA = 12'b111111010110;
            14'b11_101101111111: DATA = 12'b111111010111;
            14'b11_101110000000: DATA = 12'b111111010111;
            14'b11_101110000001: DATA = 12'b111111011000;
            14'b11_101110000010: DATA = 12'b111111011000;
            14'b11_101110000011: DATA = 12'b111111011001;
            14'b11_101110000100: DATA = 12'b111111011010;
            14'b11_101110000101: DATA = 12'b111111011010;
            14'b11_101110000110: DATA = 12'b111111011011;
            14'b11_101110000111: DATA = 12'b111111011011;
            14'b11_101110001000: DATA = 12'b111111011100;
            14'b11_101110001001: DATA = 12'b111111011100;
            14'b11_101110001010: DATA = 12'b111111011101;
            14'b11_101110001011: DATA = 12'b111111011110;
            14'b11_101110001100: DATA = 12'b111111011110;
            14'b11_101110001101: DATA = 12'b111111011111;
            14'b11_101110001110: DATA = 12'b111111011111;
            14'b11_101110001111: DATA = 12'b111111100000;
            14'b11_101110010000: DATA = 12'b111111100000;
            14'b11_101110010001: DATA = 12'b111111100001;
            14'b11_101110010010: DATA = 12'b111111100001;
            14'b11_101110010011: DATA = 12'b111111100010;
            14'b11_101110010100: DATA = 12'b111111100010;
            14'b11_101110010101: DATA = 12'b111111100011;
            14'b11_101110010110: DATA = 12'b111111100011;
            14'b11_101110010111: DATA = 12'b111111100100;
            14'b11_101110011000: DATA = 12'b111111100101;
            14'b11_101110011001: DATA = 12'b111111100101;
            14'b11_101110011010: DATA = 12'b111111100101;
            14'b11_101110011011: DATA = 12'b111111100110;
            14'b11_101110011100: DATA = 12'b111111100110;
            14'b11_101110011101: DATA = 12'b111111100111;
            14'b11_101110011110: DATA = 12'b111111100111;
            14'b11_101110011111: DATA = 12'b111111101000;
            14'b11_101110100000: DATA = 12'b111111101000;
            14'b11_101110100001: DATA = 12'b111111101001;
            14'b11_101110100010: DATA = 12'b111111101001;
            14'b11_101110100011: DATA = 12'b111111101010;
            14'b11_101110100100: DATA = 12'b111111101010;
            14'b11_101110100101: DATA = 12'b111111101011;
            14'b11_101110100110: DATA = 12'b111111101011;
            14'b11_101110100111: DATA = 12'b111111101011;
            14'b11_101110101000: DATA = 12'b111111101100;
            14'b11_101110101001: DATA = 12'b111111101100;
            14'b11_101110101010: DATA = 12'b111111101101;
            14'b11_101110101011: DATA = 12'b111111101101;
            14'b11_101110101100: DATA = 12'b111111101110;
            14'b11_101110101101: DATA = 12'b111111101110;
            14'b11_101110101110: DATA = 12'b111111101110;
            14'b11_101110101111: DATA = 12'b111111101111;
            14'b11_101110110000: DATA = 12'b111111101111;
            14'b11_101110110001: DATA = 12'b111111101111;
            14'b11_101110110010: DATA = 12'b111111110000;
            14'b11_101110110011: DATA = 12'b111111110000;
            14'b11_101110110100: DATA = 12'b111111110001;
            14'b11_101110110101: DATA = 12'b111111110001;
            14'b11_101110110110: DATA = 12'b111111110001;
            14'b11_101110110111: DATA = 12'b111111110010;
            14'b11_101110111000: DATA = 12'b111111110010;
            14'b11_101110111001: DATA = 12'b111111110010;
            14'b11_101110111010: DATA = 12'b111111110011;
            14'b11_101110111011: DATA = 12'b111111110011;
            14'b11_101110111100: DATA = 12'b111111110011;
            14'b11_101110111101: DATA = 12'b111111110100;
            14'b11_101110111110: DATA = 12'b111111110100;
            14'b11_101110111111: DATA = 12'b111111110100;
            14'b11_101111000000: DATA = 12'b111111110101;
            14'b11_101111000001: DATA = 12'b111111110101;
            14'b11_101111000010: DATA = 12'b111111110101;
            14'b11_101111000011: DATA = 12'b111111110110;
            14'b11_101111000100: DATA = 12'b111111110110;
            14'b11_101111000101: DATA = 12'b111111110110;
            14'b11_101111000110: DATA = 12'b111111110110;
            14'b11_101111000111: DATA = 12'b111111110111;
            14'b11_101111001000: DATA = 12'b111111110111;
            14'b11_101111001001: DATA = 12'b111111110111;
            14'b11_101111001010: DATA = 12'b111111110111;
            14'b11_101111001011: DATA = 12'b111111111000;
            14'b11_101111001100: DATA = 12'b111111111000;
            14'b11_101111001101: DATA = 12'b111111111000;
            14'b11_101111001110: DATA = 12'b111111111000;
            14'b11_101111001111: DATA = 12'b111111111001;
            14'b11_101111010000: DATA = 12'b111111111001;
            14'b11_101111010001: DATA = 12'b111111111001;
            14'b11_101111010010: DATA = 12'b111111111001;
            14'b11_101111010011: DATA = 12'b111111111010;
            14'b11_101111010100: DATA = 12'b111111111010;
            14'b11_101111010101: DATA = 12'b111111111010;
            14'b11_101111010110: DATA = 12'b111111111010;
            14'b11_101111010111: DATA = 12'b111111111010;
            14'b11_101111011000: DATA = 12'b111111111011;
            14'b11_101111011001: DATA = 12'b111111111011;
            14'b11_101111011010: DATA = 12'b111111111011;
            14'b11_101111011011: DATA = 12'b111111111011;
            14'b11_101111011100: DATA = 12'b111111111011;
            14'b11_101111011101: DATA = 12'b111111111100;
            14'b11_101111011110: DATA = 12'b111111111100;
            14'b11_101111011111: DATA = 12'b111111111100;
            14'b11_101111100000: DATA = 12'b111111111100;
            14'b11_101111100001: DATA = 12'b111111111100;
            14'b11_101111100010: DATA = 12'b111111111100;
            14'b11_101111100011: DATA = 12'b111111111100;
            14'b11_101111100100: DATA = 12'b111111111101;
            14'b11_101111100101: DATA = 12'b111111111101;
            14'b11_101111100110: DATA = 12'b111111111101;
            14'b11_101111100111: DATA = 12'b111111111101;
            14'b11_101111101000: DATA = 12'b111111111101;
            14'b11_101111101001: DATA = 12'b111111111101;
            14'b11_101111101010: DATA = 12'b111111111101;
            14'b11_101111101011: DATA = 12'b111111111101;
            14'b11_101111101100: DATA = 12'b111111111110;
            14'b11_101111101101: DATA = 12'b111111111110;
            14'b11_101111101110: DATA = 12'b111111111110;
            14'b11_101111101111: DATA = 12'b111111111110;
            14'b11_101111110000: DATA = 12'b111111111110;
            14'b11_101111110001: DATA = 12'b111111111110;
            14'b11_101111110010: DATA = 12'b111111111110;
            14'b11_101111110011: DATA = 12'b111111111110;
            14'b11_101111110100: DATA = 12'b111111111110;
            14'b11_101111110101: DATA = 12'b111111111110;
            14'b11_101111110110: DATA = 12'b111111111110;
            14'b11_101111110111: DATA = 12'b111111111110;
            14'b11_101111111000: DATA = 12'b111111111110;
            14'b11_101111111001: DATA = 12'b111111111110;
            14'b11_101111111010: DATA = 12'b111111111110;
            14'b11_101111111011: DATA = 12'b111111111110;
            14'b11_101111111100: DATA = 12'b111111111110;
            14'b11_101111111101: DATA = 12'b111111111110;
            14'b11_101111111110: DATA = 12'b111111111110;
            14'b11_101111111111: DATA = 12'b111111111110;
            14'b11_110000000000: DATA = 12'b111111111111;
            14'b11_110000000001: DATA = 12'b111111111110;
            14'b11_110000000010: DATA = 12'b111111111110;
            14'b11_110000000011: DATA = 12'b111111111110;
            14'b11_110000000100: DATA = 12'b111111111110;
            14'b11_110000000101: DATA = 12'b111111111110;
            14'b11_110000000110: DATA = 12'b111111111110;
            14'b11_110000000111: DATA = 12'b111111111110;
            14'b11_110000001000: DATA = 12'b111111111110;
            14'b11_110000001001: DATA = 12'b111111111110;
            14'b11_110000001010: DATA = 12'b111111111110;
            14'b11_110000001011: DATA = 12'b111111111110;
            14'b11_110000001100: DATA = 12'b111111111110;
            14'b11_110000001101: DATA = 12'b111111111110;
            14'b11_110000001110: DATA = 12'b111111111110;
            14'b11_110000001111: DATA = 12'b111111111110;
            14'b11_110000010000: DATA = 12'b111111111110;
            14'b11_110000010001: DATA = 12'b111111111110;
            14'b11_110000010010: DATA = 12'b111111111110;
            14'b11_110000010011: DATA = 12'b111111111110;
            14'b11_110000010100: DATA = 12'b111111111110;
            14'b11_110000010101: DATA = 12'b111111111101;
            14'b11_110000010110: DATA = 12'b111111111101;
            14'b11_110000010111: DATA = 12'b111111111101;
            14'b11_110000011000: DATA = 12'b111111111101;
            14'b11_110000011001: DATA = 12'b111111111101;
            14'b11_110000011010: DATA = 12'b111111111101;
            14'b11_110000011011: DATA = 12'b111111111101;
            14'b11_110000011100: DATA = 12'b111111111101;
            14'b11_110000011101: DATA = 12'b111111111100;
            14'b11_110000011110: DATA = 12'b111111111100;
            14'b11_110000011111: DATA = 12'b111111111100;
            14'b11_110000100000: DATA = 12'b111111111100;
            14'b11_110000100001: DATA = 12'b111111111100;
            14'b11_110000100010: DATA = 12'b111111111100;
            14'b11_110000100011: DATA = 12'b111111111100;
            14'b11_110000100100: DATA = 12'b111111111011;
            14'b11_110000100101: DATA = 12'b111111111011;
            14'b11_110000100110: DATA = 12'b111111111011;
            14'b11_110000100111: DATA = 12'b111111111011;
            14'b11_110000101000: DATA = 12'b111111111011;
            14'b11_110000101001: DATA = 12'b111111111010;
            14'b11_110000101010: DATA = 12'b111111111010;
            14'b11_110000101011: DATA = 12'b111111111010;
            14'b11_110000101100: DATA = 12'b111111111010;
            14'b11_110000101101: DATA = 12'b111111111010;
            14'b11_110000101110: DATA = 12'b111111111001;
            14'b11_110000101111: DATA = 12'b111111111001;
            14'b11_110000110000: DATA = 12'b111111111001;
            14'b11_110000110001: DATA = 12'b111111111001;
            14'b11_110000110010: DATA = 12'b111111111000;
            14'b11_110000110011: DATA = 12'b111111111000;
            14'b11_110000110100: DATA = 12'b111111111000;
            14'b11_110000110101: DATA = 12'b111111111000;
            14'b11_110000110110: DATA = 12'b111111110111;
            14'b11_110000110111: DATA = 12'b111111110111;
            14'b11_110000111000: DATA = 12'b111111110111;
            14'b11_110000111001: DATA = 12'b111111110111;
            14'b11_110000111010: DATA = 12'b111111110110;
            14'b11_110000111011: DATA = 12'b111111110110;
            14'b11_110000111100: DATA = 12'b111111110110;
            14'b11_110000111101: DATA = 12'b111111110110;
            14'b11_110000111110: DATA = 12'b111111110101;
            14'b11_110000111111: DATA = 12'b111111110101;
            14'b11_110001000000: DATA = 12'b111111110101;
            14'b11_110001000001: DATA = 12'b111111110100;
            14'b11_110001000010: DATA = 12'b111111110100;
            14'b11_110001000011: DATA = 12'b111111110100;
            14'b11_110001000100: DATA = 12'b111111110011;
            14'b11_110001000101: DATA = 12'b111111110011;
            14'b11_110001000110: DATA = 12'b111111110011;
            14'b11_110001000111: DATA = 12'b111111110010;
            14'b11_110001001000: DATA = 12'b111111110010;
            14'b11_110001001001: DATA = 12'b111111110010;
            14'b11_110001001010: DATA = 12'b111111110001;
            14'b11_110001001011: DATA = 12'b111111110001;
            14'b11_110001001100: DATA = 12'b111111110001;
            14'b11_110001001101: DATA = 12'b111111110000;
            14'b11_110001001110: DATA = 12'b111111110000;
            14'b11_110001001111: DATA = 12'b111111101111;
            14'b11_110001010000: DATA = 12'b111111101111;
            14'b11_110001010001: DATA = 12'b111111101111;
            14'b11_110001010010: DATA = 12'b111111101110;
            14'b11_110001010011: DATA = 12'b111111101110;
            14'b11_110001010100: DATA = 12'b111111101110;
            14'b11_110001010101: DATA = 12'b111111101101;
            14'b11_110001010110: DATA = 12'b111111101101;
            14'b11_110001010111: DATA = 12'b111111101100;
            14'b11_110001011000: DATA = 12'b111111101100;
            14'b11_110001011001: DATA = 12'b111111101011;
            14'b11_110001011010: DATA = 12'b111111101011;
            14'b11_110001011011: DATA = 12'b111111101011;
            14'b11_110001011100: DATA = 12'b111111101010;
            14'b11_110001011101: DATA = 12'b111111101010;
            14'b11_110001011110: DATA = 12'b111111101001;
            14'b11_110001011111: DATA = 12'b111111101001;
            14'b11_110001100000: DATA = 12'b111111101000;
            14'b11_110001100001: DATA = 12'b111111101000;
            14'b11_110001100010: DATA = 12'b111111100111;
            14'b11_110001100011: DATA = 12'b111111100111;
            14'b11_110001100100: DATA = 12'b111111100110;
            14'b11_110001100101: DATA = 12'b111111100110;
            14'b11_110001100110: DATA = 12'b111111100101;
            14'b11_110001100111: DATA = 12'b111111100101;
            14'b11_110001101000: DATA = 12'b111111100101;
            14'b11_110001101001: DATA = 12'b111111100100;
            14'b11_110001101010: DATA = 12'b111111100011;
            14'b11_110001101011: DATA = 12'b111111100011;
            14'b11_110001101100: DATA = 12'b111111100010;
            14'b11_110001101101: DATA = 12'b111111100010;
            14'b11_110001101110: DATA = 12'b111111100001;
            14'b11_110001101111: DATA = 12'b111111100001;
            14'b11_110001110000: DATA = 12'b111111100000;
            14'b11_110001110001: DATA = 12'b111111100000;
            14'b11_110001110010: DATA = 12'b111111011111;
            14'b11_110001110011: DATA = 12'b111111011111;
            14'b11_110001110100: DATA = 12'b111111011110;
            14'b11_110001110101: DATA = 12'b111111011110;
            14'b11_110001110110: DATA = 12'b111111011101;
            14'b11_110001110111: DATA = 12'b111111011100;
            14'b11_110001111000: DATA = 12'b111111011100;
            14'b11_110001111001: DATA = 12'b111111011011;
            14'b11_110001111010: DATA = 12'b111111011011;
            14'b11_110001111011: DATA = 12'b111111011010;
            14'b11_110001111100: DATA = 12'b111111011010;
            14'b11_110001111101: DATA = 12'b111111011001;
            14'b11_110001111110: DATA = 12'b111111011000;
            14'b11_110001111111: DATA = 12'b111111011000;
            14'b11_110010000000: DATA = 12'b111111010111;
            14'b11_110010000001: DATA = 12'b111111010111;
            14'b11_110010000010: DATA = 12'b111111010110;
            14'b11_110010000011: DATA = 12'b111111010101;
            14'b11_110010000100: DATA = 12'b111111010101;
            14'b11_110010000101: DATA = 12'b111111010100;
            14'b11_110010000110: DATA = 12'b111111010011;
            14'b11_110010000111: DATA = 12'b111111010011;
            14'b11_110010001000: DATA = 12'b111111010010;
            14'b11_110010001001: DATA = 12'b111111010001;
            14'b11_110010001010: DATA = 12'b111111010001;
            14'b11_110010001011: DATA = 12'b111111010000;
            14'b11_110010001100: DATA = 12'b111111001111;
            14'b11_110010001101: DATA = 12'b111111001111;
            14'b11_110010001110: DATA = 12'b111111001110;
            14'b11_110010001111: DATA = 12'b111111001101;
            14'b11_110010010000: DATA = 12'b111111001101;
            14'b11_110010010001: DATA = 12'b111111001100;
            14'b11_110010010010: DATA = 12'b111111001011;
            14'b11_110010010011: DATA = 12'b111111001011;
            14'b11_110010010100: DATA = 12'b111111001010;
            14'b11_110010010101: DATA = 12'b111111001001;
            14'b11_110010010110: DATA = 12'b111111001001;
            14'b11_110010010111: DATA = 12'b111111001000;
            14'b11_110010011000: DATA = 12'b111111000111;
            14'b11_110010011001: DATA = 12'b111111000110;
            14'b11_110010011010: DATA = 12'b111111000110;
            14'b11_110010011011: DATA = 12'b111111000101;
            14'b11_110010011100: DATA = 12'b111111000100;
            14'b11_110010011101: DATA = 12'b111111000011;
            14'b11_110010011110: DATA = 12'b111111000011;
            14'b11_110010011111: DATA = 12'b111111000010;
            14'b11_110010100000: DATA = 12'b111111000001;
            14'b11_110010100001: DATA = 12'b111111000000;
            14'b11_110010100010: DATA = 12'b111111000000;
            14'b11_110010100011: DATA = 12'b111110111111;
            14'b11_110010100100: DATA = 12'b111110111110;
            14'b11_110010100101: DATA = 12'b111110111101;
            14'b11_110010100110: DATA = 12'b111110111100;
            14'b11_110010100111: DATA = 12'b111110111100;
            14'b11_110010101000: DATA = 12'b111110111011;
            14'b11_110010101001: DATA = 12'b111110111010;
            14'b11_110010101010: DATA = 12'b111110111001;
            14'b11_110010101011: DATA = 12'b111110111000;
            14'b11_110010101100: DATA = 12'b111110111000;
            14'b11_110010101101: DATA = 12'b111110110111;
            14'b11_110010101110: DATA = 12'b111110110110;
            14'b11_110010101111: DATA = 12'b111110110101;
            14'b11_110010110000: DATA = 12'b111110110100;
            14'b11_110010110001: DATA = 12'b111110110100;
            14'b11_110010110010: DATA = 12'b111110110011;
            14'b11_110010110011: DATA = 12'b111110110010;
            14'b11_110010110100: DATA = 12'b111110110001;
            14'b11_110010110101: DATA = 12'b111110110000;
            14'b11_110010110110: DATA = 12'b111110101111;
            14'b11_110010110111: DATA = 12'b111110101110;
            14'b11_110010111000: DATA = 12'b111110101110;
            14'b11_110010111001: DATA = 12'b111110101101;
            14'b11_110010111010: DATA = 12'b111110101100;
            14'b11_110010111011: DATA = 12'b111110101011;
            14'b11_110010111100: DATA = 12'b111110101010;
            14'b11_110010111101: DATA = 12'b111110101001;
            14'b11_110010111110: DATA = 12'b111110101000;
            14'b11_110010111111: DATA = 12'b111110100111;
            14'b11_110011000000: DATA = 12'b111110100110;
            14'b11_110011000001: DATA = 12'b111110100101;
            14'b11_110011000010: DATA = 12'b111110100101;
            14'b11_110011000011: DATA = 12'b111110100100;
            14'b11_110011000100: DATA = 12'b111110100011;
            14'b11_110011000101: DATA = 12'b111110100010;
            14'b11_110011000110: DATA = 12'b111110100001;
            14'b11_110011000111: DATA = 12'b111110100000;
            14'b11_110011001000: DATA = 12'b111110011111;
            14'b11_110011001001: DATA = 12'b111110011110;
            14'b11_110011001010: DATA = 12'b111110011101;
            14'b11_110011001011: DATA = 12'b111110011100;
            14'b11_110011001100: DATA = 12'b111110011011;
            14'b11_110011001101: DATA = 12'b111110011010;
            14'b11_110011001110: DATA = 12'b111110011001;
            14'b11_110011001111: DATA = 12'b111110011000;
            14'b11_110011010000: DATA = 12'b111110010111;
            14'b11_110011010001: DATA = 12'b111110010110;
            14'b11_110011010010: DATA = 12'b111110010101;
            14'b11_110011010011: DATA = 12'b111110010100;
            14'b11_110011010100: DATA = 12'b111110010011;
            14'b11_110011010101: DATA = 12'b111110010010;
            14'b11_110011010110: DATA = 12'b111110010001;
            14'b11_110011010111: DATA = 12'b111110010000;
            14'b11_110011011000: DATA = 12'b111110001111;
            14'b11_110011011001: DATA = 12'b111110001110;
            14'b11_110011011010: DATA = 12'b111110001101;
            14'b11_110011011011: DATA = 12'b111110001100;
            14'b11_110011011100: DATA = 12'b111110001011;
            14'b11_110011011101: DATA = 12'b111110001010;
            14'b11_110011011110: DATA = 12'b111110001001;
            14'b11_110011011111: DATA = 12'b111110001000;
            14'b11_110011100000: DATA = 12'b111110000111;
            14'b11_110011100001: DATA = 12'b111110000110;
            14'b11_110011100010: DATA = 12'b111110000101;
            14'b11_110011100011: DATA = 12'b111110000100;
            14'b11_110011100100: DATA = 12'b111110000011;
            14'b11_110011100101: DATA = 12'b111110000001;
            14'b11_110011100110: DATA = 12'b111110000000;
            14'b11_110011100111: DATA = 12'b111101111111;
            14'b11_110011101000: DATA = 12'b111101111110;
            14'b11_110011101001: DATA = 12'b111101111101;
            14'b11_110011101010: DATA = 12'b111101111100;
            14'b11_110011101011: DATA = 12'b111101111011;
            14'b11_110011101100: DATA = 12'b111101111010;
            14'b11_110011101101: DATA = 12'b111101111001;
            14'b11_110011101110: DATA = 12'b111101111000;
            14'b11_110011101111: DATA = 12'b111101110110;
            14'b11_110011110000: DATA = 12'b111101110101;
            14'b11_110011110001: DATA = 12'b111101110100;
            14'b11_110011110010: DATA = 12'b111101110011;
            14'b11_110011110011: DATA = 12'b111101110010;
            14'b11_110011110100: DATA = 12'b111101110001;
            14'b11_110011110101: DATA = 12'b111101110000;
            14'b11_110011110110: DATA = 12'b111101101110;
            14'b11_110011110111: DATA = 12'b111101101101;
            14'b11_110011111000: DATA = 12'b111101101100;
            14'b11_110011111001: DATA = 12'b111101101011;
            14'b11_110011111010: DATA = 12'b111101101010;
            14'b11_110011111011: DATA = 12'b111101101001;
            14'b11_110011111100: DATA = 12'b111101100111;
            14'b11_110011111101: DATA = 12'b111101100110;
            14'b11_110011111110: DATA = 12'b111101100101;
            14'b11_110011111111: DATA = 12'b111101100100;
            14'b11_110100000000: DATA = 12'b111101100011;
            14'b11_110100000001: DATA = 12'b111101100001;
            14'b11_110100000010: DATA = 12'b111101100000;
            14'b11_110100000011: DATA = 12'b111101011111;
            14'b11_110100000100: DATA = 12'b111101011110;
            14'b11_110100000101: DATA = 12'b111101011101;
            14'b11_110100000110: DATA = 12'b111101011011;
            14'b11_110100000111: DATA = 12'b111101011010;
            14'b11_110100001000: DATA = 12'b111101011001;
            14'b11_110100001001: DATA = 12'b111101011000;
            14'b11_110100001010: DATA = 12'b111101010110;
            14'b11_110100001011: DATA = 12'b111101010101;
            14'b11_110100001100: DATA = 12'b111101010100;
            14'b11_110100001101: DATA = 12'b111101010011;
            14'b11_110100001110: DATA = 12'b111101010001;
            14'b11_110100001111: DATA = 12'b111101010000;
            14'b11_110100010000: DATA = 12'b111101001111;
            14'b11_110100010001: DATA = 12'b111101001110;
            14'b11_110100010010: DATA = 12'b111101001100;
            14'b11_110100010011: DATA = 12'b111101001011;
            14'b11_110100010100: DATA = 12'b111101001010;
            14'b11_110100010101: DATA = 12'b111101001000;
            14'b11_110100010110: DATA = 12'b111101000111;
            14'b11_110100010111: DATA = 12'b111101000110;
            14'b11_110100011000: DATA = 12'b111101000101;
            14'b11_110100011001: DATA = 12'b111101000011;
            14'b11_110100011010: DATA = 12'b111101000010;
            14'b11_110100011011: DATA = 12'b111101000001;
            14'b11_110100011100: DATA = 12'b111100111111;
            14'b11_110100011101: DATA = 12'b111100111110;
            14'b11_110100011110: DATA = 12'b111100111101;
            14'b11_110100011111: DATA = 12'b111100111011;
            14'b11_110100100000: DATA = 12'b111100111010;
            14'b11_110100100001: DATA = 12'b111100111001;
            14'b11_110100100010: DATA = 12'b111100110111;
            14'b11_110100100011: DATA = 12'b111100110110;
            14'b11_110100100100: DATA = 12'b111100110101;
            14'b11_110100100101: DATA = 12'b111100110011;
            14'b11_110100100110: DATA = 12'b111100110010;
            14'b11_110100100111: DATA = 12'b111100110000;
            14'b11_110100101000: DATA = 12'b111100101111;
            14'b11_110100101001: DATA = 12'b111100101110;
            14'b11_110100101010: DATA = 12'b111100101100;
            14'b11_110100101011: DATA = 12'b111100101011;
            14'b11_110100101100: DATA = 12'b111100101010;
            14'b11_110100101101: DATA = 12'b111100101000;
            14'b11_110100101110: DATA = 12'b111100100111;
            14'b11_110100101111: DATA = 12'b111100100101;
            14'b11_110100110000: DATA = 12'b111100100100;
            14'b11_110100110001: DATA = 12'b111100100011;
            14'b11_110100110010: DATA = 12'b111100100001;
            14'b11_110100110011: DATA = 12'b111100100000;
            14'b11_110100110100: DATA = 12'b111100011110;
            14'b11_110100110101: DATA = 12'b111100011101;
            14'b11_110100110110: DATA = 12'b111100011011;
            14'b11_110100110111: DATA = 12'b111100011010;
            14'b11_110100111000: DATA = 12'b111100011000;
            14'b11_110100111001: DATA = 12'b111100010111;
            14'b11_110100111010: DATA = 12'b111100010110;
            14'b11_110100111011: DATA = 12'b111100010100;
            14'b11_110100111100: DATA = 12'b111100010011;
            14'b11_110100111101: DATA = 12'b111100010001;
            14'b11_110100111110: DATA = 12'b111100010000;
            14'b11_110100111111: DATA = 12'b111100001110;
            14'b11_110101000000: DATA = 12'b111100001101;
            14'b11_110101000001: DATA = 12'b111100001011;
            14'b11_110101000010: DATA = 12'b111100001010;
            14'b11_110101000011: DATA = 12'b111100001000;
            14'b11_110101000100: DATA = 12'b111100000111;
            14'b11_110101000101: DATA = 12'b111100000101;
            14'b11_110101000110: DATA = 12'b111100000100;
            14'b11_110101000111: DATA = 12'b111100000010;
            14'b11_110101001000: DATA = 12'b111100000001;
            14'b11_110101001001: DATA = 12'b111011111111;
            14'b11_110101001010: DATA = 12'b111011111110;
            14'b11_110101001011: DATA = 12'b111011111100;
            14'b11_110101001100: DATA = 12'b111011111011;
            14'b11_110101001101: DATA = 12'b111011111001;
            14'b11_110101001110: DATA = 12'b111011111000;
            14'b11_110101001111: DATA = 12'b111011110110;
            14'b11_110101010000: DATA = 12'b111011110101;
            14'b11_110101010001: DATA = 12'b111011110011;
            14'b11_110101010010: DATA = 12'b111011110001;
            14'b11_110101010011: DATA = 12'b111011110000;
            14'b11_110101010100: DATA = 12'b111011101110;
            14'b11_110101010101: DATA = 12'b111011101101;
            14'b11_110101010110: DATA = 12'b111011101011;
            14'b11_110101010111: DATA = 12'b111011101010;
            14'b11_110101011000: DATA = 12'b111011101000;
            14'b11_110101011001: DATA = 12'b111011100110;
            14'b11_110101011010: DATA = 12'b111011100101;
            14'b11_110101011011: DATA = 12'b111011100011;
            14'b11_110101011100: DATA = 12'b111011100010;
            14'b11_110101011101: DATA = 12'b111011100000;
            14'b11_110101011110: DATA = 12'b111011011110;
            14'b11_110101011111: DATA = 12'b111011011101;
            14'b11_110101100000: DATA = 12'b111011011011;
            14'b11_110101100001: DATA = 12'b111011011010;
            14'b11_110101100010: DATA = 12'b111011011000;
            14'b11_110101100011: DATA = 12'b111011010110;
            14'b11_110101100100: DATA = 12'b111011010101;
            14'b11_110101100101: DATA = 12'b111011010011;
            14'b11_110101100110: DATA = 12'b111011010010;
            14'b11_110101100111: DATA = 12'b111011010000;
            14'b11_110101101000: DATA = 12'b111011001110;
            14'b11_110101101001: DATA = 12'b111011001101;
            14'b11_110101101010: DATA = 12'b111011001011;
            14'b11_110101101011: DATA = 12'b111011001001;
            14'b11_110101101100: DATA = 12'b111011001000;
            14'b11_110101101101: DATA = 12'b111011000110;
            14'b11_110101101110: DATA = 12'b111011000100;
            14'b11_110101101111: DATA = 12'b111011000011;
            14'b11_110101110000: DATA = 12'b111011000001;
            14'b11_110101110001: DATA = 12'b111010111111;
            14'b11_110101110010: DATA = 12'b111010111110;
            14'b11_110101110011: DATA = 12'b111010111100;
            14'b11_110101110100: DATA = 12'b111010111010;
            14'b11_110101110101: DATA = 12'b111010111000;
            14'b11_110101110110: DATA = 12'b111010110111;
            14'b11_110101110111: DATA = 12'b111010110101;
            14'b11_110101111000: DATA = 12'b111010110011;
            14'b11_110101111001: DATA = 12'b111010110010;
            14'b11_110101111010: DATA = 12'b111010110000;
            14'b11_110101111011: DATA = 12'b111010101110;
            14'b11_110101111100: DATA = 12'b111010101100;
            14'b11_110101111101: DATA = 12'b111010101011;
            14'b11_110101111110: DATA = 12'b111010101001;
            14'b11_110101111111: DATA = 12'b111010100111;
            14'b11_110110000000: DATA = 12'b111010100110;
            14'b11_110110000001: DATA = 12'b111010100100;
            14'b11_110110000010: DATA = 12'b111010100010;
            14'b11_110110000011: DATA = 12'b111010100000;
            14'b11_110110000100: DATA = 12'b111010011111;
            14'b11_110110000101: DATA = 12'b111010011101;
            14'b11_110110000110: DATA = 12'b111010011011;
            14'b11_110110000111: DATA = 12'b111010011001;
            14'b11_110110001000: DATA = 12'b111010010111;
            14'b11_110110001001: DATA = 12'b111010010110;
            14'b11_110110001010: DATA = 12'b111010010100;
            14'b11_110110001011: DATA = 12'b111010010010;
            14'b11_110110001100: DATA = 12'b111010010000;
            14'b11_110110001101: DATA = 12'b111010001111;
            14'b11_110110001110: DATA = 12'b111010001101;
            14'b11_110110001111: DATA = 12'b111010001011;
            14'b11_110110010000: DATA = 12'b111010001001;
            14'b11_110110010001: DATA = 12'b111010000111;
            14'b11_110110010010: DATA = 12'b111010000101;
            14'b11_110110010011: DATA = 12'b111010000100;
            14'b11_110110010100: DATA = 12'b111010000010;
            14'b11_110110010101: DATA = 12'b111010000000;
            14'b11_110110010110: DATA = 12'b111001111110;
            14'b11_110110010111: DATA = 12'b111001111100;
            14'b11_110110011000: DATA = 12'b111001111011;
            14'b11_110110011001: DATA = 12'b111001111001;
            14'b11_110110011010: DATA = 12'b111001110111;
            14'b11_110110011011: DATA = 12'b111001110101;
            14'b11_110110011100: DATA = 12'b111001110011;
            14'b11_110110011101: DATA = 12'b111001110001;
            14'b11_110110011110: DATA = 12'b111001101111;
            14'b11_110110011111: DATA = 12'b111001101110;
            14'b11_110110100000: DATA = 12'b111001101100;
            14'b11_110110100001: DATA = 12'b111001101010;
            14'b11_110110100010: DATA = 12'b111001101000;
            14'b11_110110100011: DATA = 12'b111001100110;
            14'b11_110110100100: DATA = 12'b111001100100;
            14'b11_110110100101: DATA = 12'b111001100010;
            14'b11_110110100110: DATA = 12'b111001100000;
            14'b11_110110100111: DATA = 12'b111001011110;
            14'b11_110110101000: DATA = 12'b111001011101;
            14'b11_110110101001: DATA = 12'b111001011011;
            14'b11_110110101010: DATA = 12'b111001011001;
            14'b11_110110101011: DATA = 12'b111001010111;
            14'b11_110110101100: DATA = 12'b111001010101;
            14'b11_110110101101: DATA = 12'b111001010011;
            14'b11_110110101110: DATA = 12'b111001010001;
            14'b11_110110101111: DATA = 12'b111001001111;
            14'b11_110110110000: DATA = 12'b111001001101;
            14'b11_110110110001: DATA = 12'b111001001011;
            14'b11_110110110010: DATA = 12'b111001001001;
            14'b11_110110110011: DATA = 12'b111001000111;
            14'b11_110110110100: DATA = 12'b111001000101;
            14'b11_110110110101: DATA = 12'b111001000100;
            14'b11_110110110110: DATA = 12'b111001000010;
            14'b11_110110110111: DATA = 12'b111001000000;
            14'b11_110110111000: DATA = 12'b111000111110;
            14'b11_110110111001: DATA = 12'b111000111100;
            14'b11_110110111010: DATA = 12'b111000111010;
            14'b11_110110111011: DATA = 12'b111000111000;
            14'b11_110110111100: DATA = 12'b111000110110;
            14'b11_110110111101: DATA = 12'b111000110100;
            14'b11_110110111110: DATA = 12'b111000110010;
            14'b11_110110111111: DATA = 12'b111000110000;
            14'b11_110111000000: DATA = 12'b111000101110;
            14'b11_110111000001: DATA = 12'b111000101100;
            14'b11_110111000010: DATA = 12'b111000101010;
            14'b11_110111000011: DATA = 12'b111000101000;
            14'b11_110111000100: DATA = 12'b111000100110;
            14'b11_110111000101: DATA = 12'b111000100100;
            14'b11_110111000110: DATA = 12'b111000100010;
            14'b11_110111000111: DATA = 12'b111000100000;
            14'b11_110111001000: DATA = 12'b111000011110;
            14'b11_110111001001: DATA = 12'b111000011100;
            14'b11_110111001010: DATA = 12'b111000011010;
            14'b11_110111001011: DATA = 12'b111000011000;
            14'b11_110111001100: DATA = 12'b111000010110;
            14'b11_110111001101: DATA = 12'b111000010100;
            14'b11_110111001110: DATA = 12'b111000010010;
            14'b11_110111001111: DATA = 12'b111000010000;
            14'b11_110111010000: DATA = 12'b111000001110;
            14'b11_110111010001: DATA = 12'b111000001011;
            14'b11_110111010010: DATA = 12'b111000001001;
            14'b11_110111010011: DATA = 12'b111000000111;
            14'b11_110111010100: DATA = 12'b111000000101;
            14'b11_110111010101: DATA = 12'b111000000011;
            14'b11_110111010110: DATA = 12'b111000000001;
            14'b11_110111010111: DATA = 12'b110111111111;
            14'b11_110111011000: DATA = 12'b110111111101;
            14'b11_110111011001: DATA = 12'b110111111011;
            14'b11_110111011010: DATA = 12'b110111111001;
            14'b11_110111011011: DATA = 12'b110111110111;
            14'b11_110111011100: DATA = 12'b110111110101;
            14'b11_110111011101: DATA = 12'b110111110011;
            14'b11_110111011110: DATA = 12'b110111110000;
            14'b11_110111011111: DATA = 12'b110111101110;
            14'b11_110111100000: DATA = 12'b110111101100;
            14'b11_110111100001: DATA = 12'b110111101010;
            14'b11_110111100010: DATA = 12'b110111101000;
            14'b11_110111100011: DATA = 12'b110111100110;
            14'b11_110111100100: DATA = 12'b110111100100;
            14'b11_110111100101: DATA = 12'b110111100010;
            14'b11_110111100110: DATA = 12'b110111100000;
            14'b11_110111100111: DATA = 12'b110111011101;
            14'b11_110111101000: DATA = 12'b110111011011;
            14'b11_110111101001: DATA = 12'b110111011001;
            14'b11_110111101010: DATA = 12'b110111010111;
            14'b11_110111101011: DATA = 12'b110111010101;
            14'b11_110111101100: DATA = 12'b110111010011;
            14'b11_110111101101: DATA = 12'b110111010001;
            14'b11_110111101110: DATA = 12'b110111001110;
            14'b11_110111101111: DATA = 12'b110111001100;
            14'b11_110111110000: DATA = 12'b110111001010;
            14'b11_110111110001: DATA = 12'b110111001000;
            14'b11_110111110010: DATA = 12'b110111000110;
            14'b11_110111110011: DATA = 12'b110111000100;
            14'b11_110111110100: DATA = 12'b110111000001;
            14'b11_110111110101: DATA = 12'b110110111111;
            14'b11_110111110110: DATA = 12'b110110111101;
            14'b11_110111110111: DATA = 12'b110110111011;
            14'b11_110111111000: DATA = 12'b110110111001;
            14'b11_110111111001: DATA = 12'b110110110110;
            14'b11_110111111010: DATA = 12'b110110110100;
            14'b11_110111111011: DATA = 12'b110110110010;
            14'b11_110111111100: DATA = 12'b110110110000;
            14'b11_110111111101: DATA = 12'b110110101110;
            14'b11_110111111110: DATA = 12'b110110101011;
            14'b11_110111111111: DATA = 12'b110110101001;
            14'b11_111000000000: DATA = 12'b110110100111;
            14'b11_111000000001: DATA = 12'b110110100101;
            14'b11_111000000010: DATA = 12'b110110100011;
            14'b11_111000000011: DATA = 12'b110110100000;
            14'b11_111000000100: DATA = 12'b110110011110;
            14'b11_111000000101: DATA = 12'b110110011100;
            14'b11_111000000110: DATA = 12'b110110011010;
            14'b11_111000000111: DATA = 12'b110110010111;
            14'b11_111000001000: DATA = 12'b110110010101;
            14'b11_111000001001: DATA = 12'b110110010011;
            14'b11_111000001010: DATA = 12'b110110010001;
            14'b11_111000001011: DATA = 12'b110110001110;
            14'b11_111000001100: DATA = 12'b110110001100;
            14'b11_111000001101: DATA = 12'b110110001010;
            14'b11_111000001110: DATA = 12'b110110001000;
            14'b11_111000001111: DATA = 12'b110110000101;
            14'b11_111000010000: DATA = 12'b110110000011;
            14'b11_111000010001: DATA = 12'b110110000001;
            14'b11_111000010010: DATA = 12'b110101111110;
            14'b11_111000010011: DATA = 12'b110101111100;
            14'b11_111000010100: DATA = 12'b110101111010;
            14'b11_111000010101: DATA = 12'b110101111000;
            14'b11_111000010110: DATA = 12'b110101110101;
            14'b11_111000010111: DATA = 12'b110101110011;
            14'b11_111000011000: DATA = 12'b110101110001;
            14'b11_111000011001: DATA = 12'b110101101110;
            14'b11_111000011010: DATA = 12'b110101101100;
            14'b11_111000011011: DATA = 12'b110101101010;
            14'b11_111000011100: DATA = 12'b110101100111;
            14'b11_111000011101: DATA = 12'b110101100101;
            14'b11_111000011110: DATA = 12'b110101100011;
            14'b11_111000011111: DATA = 12'b110101100001;
            14'b11_111000100000: DATA = 12'b110101011110;
            14'b11_111000100001: DATA = 12'b110101011100;
            14'b11_111000100010: DATA = 12'b110101011010;
            14'b11_111000100011: DATA = 12'b110101010111;
            14'b11_111000100100: DATA = 12'b110101010101;
            14'b11_111000100101: DATA = 12'b110101010011;
            14'b11_111000100110: DATA = 12'b110101010000;
            14'b11_111000100111: DATA = 12'b110101001110;
            14'b11_111000101000: DATA = 12'b110101001011;
            14'b11_111000101001: DATA = 12'b110101001001;
            14'b11_111000101010: DATA = 12'b110101000111;
            14'b11_111000101011: DATA = 12'b110101000100;
            14'b11_111000101100: DATA = 12'b110101000010;
            14'b11_111000101101: DATA = 12'b110101000000;
            14'b11_111000101110: DATA = 12'b110100111101;
            14'b11_111000101111: DATA = 12'b110100111011;
            14'b11_111000110000: DATA = 12'b110100111001;
            14'b11_111000110001: DATA = 12'b110100110110;
            14'b11_111000110010: DATA = 12'b110100110100;
            14'b11_111000110011: DATA = 12'b110100110001;
            14'b11_111000110100: DATA = 12'b110100101111;
            14'b11_111000110101: DATA = 12'b110100101101;
            14'b11_111000110110: DATA = 12'b110100101010;
            14'b11_111000110111: DATA = 12'b110100101000;
            14'b11_111000111000: DATA = 12'b110100100101;
            14'b11_111000111001: DATA = 12'b110100100011;
            14'b11_111000111010: DATA = 12'b110100100001;
            14'b11_111000111011: DATA = 12'b110100011110;
            14'b11_111000111100: DATA = 12'b110100011100;
            14'b11_111000111101: DATA = 12'b110100011001;
            14'b11_111000111110: DATA = 12'b110100010111;
            14'b11_111000111111: DATA = 12'b110100010101;
            14'b11_111001000000: DATA = 12'b110100010010;
            14'b11_111001000001: DATA = 12'b110100010000;
            14'b11_111001000010: DATA = 12'b110100001101;
            14'b11_111001000011: DATA = 12'b110100001011;
            14'b11_111001000100: DATA = 12'b110100001000;
            14'b11_111001000101: DATA = 12'b110100000110;
            14'b11_111001000110: DATA = 12'b110100000011;
            14'b11_111001000111: DATA = 12'b110100000001;
            14'b11_111001001000: DATA = 12'b110011111111;
            14'b11_111001001001: DATA = 12'b110011111100;
            14'b11_111001001010: DATA = 12'b110011111010;
            14'b11_111001001011: DATA = 12'b110011110111;
            14'b11_111001001100: DATA = 12'b110011110101;
            14'b11_111001001101: DATA = 12'b110011110010;
            14'b11_111001001110: DATA = 12'b110011110000;
            14'b11_111001001111: DATA = 12'b110011101101;
            14'b11_111001010000: DATA = 12'b110011101011;
            14'b11_111001010001: DATA = 12'b110011101000;
            14'b11_111001010010: DATA = 12'b110011100110;
            14'b11_111001010011: DATA = 12'b110011100011;
            14'b11_111001010100: DATA = 12'b110011100001;
            14'b11_111001010101: DATA = 12'b110011011110;
            14'b11_111001010110: DATA = 12'b110011011100;
            14'b11_111001010111: DATA = 12'b110011011001;
            14'b11_111001011000: DATA = 12'b110011010111;
            14'b11_111001011001: DATA = 12'b110011010100;
            14'b11_111001011010: DATA = 12'b110011010010;
            14'b11_111001011011: DATA = 12'b110011001111;
            14'b11_111001011100: DATA = 12'b110011001101;
            14'b11_111001011101: DATA = 12'b110011001010;
            14'b11_111001011110: DATA = 12'b110011001000;
            14'b11_111001011111: DATA = 12'b110011000101;
            14'b11_111001100000: DATA = 12'b110011000011;
            14'b11_111001100001: DATA = 12'b110011000000;
            14'b11_111001100010: DATA = 12'b110010111110;
            14'b11_111001100011: DATA = 12'b110010111011;
            14'b11_111001100100: DATA = 12'b110010111001;
            14'b11_111001100101: DATA = 12'b110010110110;
            14'b11_111001100110: DATA = 12'b110010110100;
            14'b11_111001100111: DATA = 12'b110010110001;
            14'b11_111001101000: DATA = 12'b110010101111;
            14'b11_111001101001: DATA = 12'b110010101100;
            14'b11_111001101010: DATA = 12'b110010101010;
            14'b11_111001101011: DATA = 12'b110010100111;
            14'b11_111001101100: DATA = 12'b110010100100;
            14'b11_111001101101: DATA = 12'b110010100010;
            14'b11_111001101110: DATA = 12'b110010011111;
            14'b11_111001101111: DATA = 12'b110010011101;
            14'b11_111001110000: DATA = 12'b110010011010;
            14'b11_111001110001: DATA = 12'b110010011000;
            14'b11_111001110010: DATA = 12'b110010010101;
            14'b11_111001110011: DATA = 12'b110010010010;
            14'b11_111001110100: DATA = 12'b110010010000;
            14'b11_111001110101: DATA = 12'b110010001101;
            14'b11_111001110110: DATA = 12'b110010001011;
            14'b11_111001110111: DATA = 12'b110010001000;
            14'b11_111001111000: DATA = 12'b110010000110;
            14'b11_111001111001: DATA = 12'b110010000011;
            14'b11_111001111010: DATA = 12'b110010000000;
            14'b11_111001111011: DATA = 12'b110001111110;
            14'b11_111001111100: DATA = 12'b110001111011;
            14'b11_111001111101: DATA = 12'b110001111001;
            14'b11_111001111110: DATA = 12'b110001110110;
            14'b11_111001111111: DATA = 12'b110001110011;
            14'b11_111010000000: DATA = 12'b110001110001;
            14'b11_111010000001: DATA = 12'b110001101110;
            14'b11_111010000010: DATA = 12'b110001101100;
            14'b11_111010000011: DATA = 12'b110001101001;
            14'b11_111010000100: DATA = 12'b110001100110;
            14'b11_111010000101: DATA = 12'b110001100100;
            14'b11_111010000110: DATA = 12'b110001100001;
            14'b11_111010000111: DATA = 12'b110001011110;
            14'b11_111010001000: DATA = 12'b110001011100;
            14'b11_111010001001: DATA = 12'b110001011001;
            14'b11_111010001010: DATA = 12'b110001010111;
            14'b11_111010001011: DATA = 12'b110001010100;
            14'b11_111010001100: DATA = 12'b110001010001;
            14'b11_111010001101: DATA = 12'b110001001111;
            14'b11_111010001110: DATA = 12'b110001001100;
            14'b11_111010001111: DATA = 12'b110001001001;
            14'b11_111010010000: DATA = 12'b110001000111;
            14'b11_111010010001: DATA = 12'b110001000100;
            14'b11_111010010010: DATA = 12'b110001000001;
            14'b11_111010010011: DATA = 12'b110000111111;
            14'b11_111010010100: DATA = 12'b110000111100;
            14'b11_111010010101: DATA = 12'b110000111001;
            14'b11_111010010110: DATA = 12'b110000110111;
            14'b11_111010010111: DATA = 12'b110000110100;
            14'b11_111010011000: DATA = 12'b110000110001;
            14'b11_111010011001: DATA = 12'b110000101111;
            14'b11_111010011010: DATA = 12'b110000101100;
            14'b11_111010011011: DATA = 12'b110000101001;
            14'b11_111010011100: DATA = 12'b110000100111;
            14'b11_111010011101: DATA = 12'b110000100100;
            14'b11_111010011110: DATA = 12'b110000100001;
            14'b11_111010011111: DATA = 12'b110000011111;
            14'b11_111010100000: DATA = 12'b110000011100;
            14'b11_111010100001: DATA = 12'b110000011001;
            14'b11_111010100010: DATA = 12'b110000010110;
            14'b11_111010100011: DATA = 12'b110000010100;
            14'b11_111010100100: DATA = 12'b110000010001;
            14'b11_111010100101: DATA = 12'b110000001110;
            14'b11_111010100110: DATA = 12'b110000001100;
            14'b11_111010100111: DATA = 12'b110000001001;
            14'b11_111010101000: DATA = 12'b110000000110;
            14'b11_111010101001: DATA = 12'b110000000100;
            14'b11_111010101010: DATA = 12'b110000000001;
            14'b11_111010101011: DATA = 12'b101111111110;
            14'b11_111010101100: DATA = 12'b101111111011;
            14'b11_111010101101: DATA = 12'b101111111001;
            14'b11_111010101110: DATA = 12'b101111110110;
            14'b11_111010101111: DATA = 12'b101111110011;
            14'b11_111010110000: DATA = 12'b101111110000;
            14'b11_111010110001: DATA = 12'b101111101110;
            14'b11_111010110010: DATA = 12'b101111101011;
            14'b11_111010110011: DATA = 12'b101111101000;
            14'b11_111010110100: DATA = 12'b101111100110;
            14'b11_111010110101: DATA = 12'b101111100011;
            14'b11_111010110110: DATA = 12'b101111100000;
            14'b11_111010110111: DATA = 12'b101111011101;
            14'b11_111010111000: DATA = 12'b101111011011;
            14'b11_111010111001: DATA = 12'b101111011000;
            14'b11_111010111010: DATA = 12'b101111010101;
            14'b11_111010111011: DATA = 12'b101111010010;
            14'b11_111010111100: DATA = 12'b101111010000;
            14'b11_111010111101: DATA = 12'b101111001101;
            14'b11_111010111110: DATA = 12'b101111001010;
            14'b11_111010111111: DATA = 12'b101111000111;
            14'b11_111011000000: DATA = 12'b101111000100;
            14'b11_111011000001: DATA = 12'b101111000010;
            14'b11_111011000010: DATA = 12'b101110111111;
            14'b11_111011000011: DATA = 12'b101110111100;
            14'b11_111011000100: DATA = 12'b101110111001;
            14'b11_111011000101: DATA = 12'b101110110111;
            14'b11_111011000110: DATA = 12'b101110110100;
            14'b11_111011000111: DATA = 12'b101110110001;
            14'b11_111011001000: DATA = 12'b101110101110;
            14'b11_111011001001: DATA = 12'b101110101011;
            14'b11_111011001010: DATA = 12'b101110101001;
            14'b11_111011001011: DATA = 12'b101110100110;
            14'b11_111011001100: DATA = 12'b101110100011;
            14'b11_111011001101: DATA = 12'b101110100000;
            14'b11_111011001110: DATA = 12'b101110011101;
            14'b11_111011001111: DATA = 12'b101110011011;
            14'b11_111011010000: DATA = 12'b101110011000;
            14'b11_111011010001: DATA = 12'b101110010101;
            14'b11_111011010010: DATA = 12'b101110010010;
            14'b11_111011010011: DATA = 12'b101110001111;
            14'b11_111011010100: DATA = 12'b101110001101;
            14'b11_111011010101: DATA = 12'b101110001010;
            14'b11_111011010110: DATA = 12'b101110000111;
            14'b11_111011010111: DATA = 12'b101110000100;
            14'b11_111011011000: DATA = 12'b101110000001;
            14'b11_111011011001: DATA = 12'b101101111111;
            14'b11_111011011010: DATA = 12'b101101111100;
            14'b11_111011011011: DATA = 12'b101101111001;
            14'b11_111011011100: DATA = 12'b101101110110;
            14'b11_111011011101: DATA = 12'b101101110011;
            14'b11_111011011110: DATA = 12'b101101110000;
            14'b11_111011011111: DATA = 12'b101101101110;
            14'b11_111011100000: DATA = 12'b101101101011;
            14'b11_111011100001: DATA = 12'b101101101000;
            14'b11_111011100010: DATA = 12'b101101100101;
            14'b11_111011100011: DATA = 12'b101101100010;
            14'b11_111011100100: DATA = 12'b101101011111;
            14'b11_111011100101: DATA = 12'b101101011100;
            14'b11_111011100110: DATA = 12'b101101011010;
            14'b11_111011100111: DATA = 12'b101101010111;
            14'b11_111011101000: DATA = 12'b101101010100;
            14'b11_111011101001: DATA = 12'b101101010001;
            14'b11_111011101010: DATA = 12'b101101001110;
            14'b11_111011101011: DATA = 12'b101101001011;
            14'b11_111011101100: DATA = 12'b101101001000;
            14'b11_111011101101: DATA = 12'b101101000110;
            14'b11_111011101110: DATA = 12'b101101000011;
            14'b11_111011101111: DATA = 12'b101101000000;
            14'b11_111011110000: DATA = 12'b101100111101;
            14'b11_111011110001: DATA = 12'b101100111010;
            14'b11_111011110010: DATA = 12'b101100110111;
            14'b11_111011110011: DATA = 12'b101100110100;
            14'b11_111011110100: DATA = 12'b101100110010;
            14'b11_111011110101: DATA = 12'b101100101111;
            14'b11_111011110110: DATA = 12'b101100101100;
            14'b11_111011110111: DATA = 12'b101100101001;
            14'b11_111011111000: DATA = 12'b101100100110;
            14'b11_111011111001: DATA = 12'b101100100011;
            14'b11_111011111010: DATA = 12'b101100100000;
            14'b11_111011111011: DATA = 12'b101100011101;
            14'b11_111011111100: DATA = 12'b101100011010;
            14'b11_111011111101: DATA = 12'b101100011000;
            14'b11_111011111110: DATA = 12'b101100010101;
            14'b11_111011111111: DATA = 12'b101100010010;
            14'b11_111100000000: DATA = 12'b101100001111;
            14'b11_111100000001: DATA = 12'b101100001100;
            14'b11_111100000010: DATA = 12'b101100001001;
            14'b11_111100000011: DATA = 12'b101100000110;
            14'b11_111100000100: DATA = 12'b101100000011;
            14'b11_111100000101: DATA = 12'b101100000000;
            14'b11_111100000110: DATA = 12'b101011111101;
            14'b11_111100000111: DATA = 12'b101011111011;
            14'b11_111100001000: DATA = 12'b101011111000;
            14'b11_111100001001: DATA = 12'b101011110101;
            14'b11_111100001010: DATA = 12'b101011110010;
            14'b11_111100001011: DATA = 12'b101011101111;
            14'b11_111100001100: DATA = 12'b101011101100;
            14'b11_111100001101: DATA = 12'b101011101001;
            14'b11_111100001110: DATA = 12'b101011100110;
            14'b11_111100001111: DATA = 12'b101011100011;
            14'b11_111100010000: DATA = 12'b101011100000;
            14'b11_111100010001: DATA = 12'b101011011101;
            14'b11_111100010010: DATA = 12'b101011011010;
            14'b11_111100010011: DATA = 12'b101011010111;
            14'b11_111100010100: DATA = 12'b101011010100;
            14'b11_111100010101: DATA = 12'b101011010010;
            14'b11_111100010110: DATA = 12'b101011001111;
            14'b11_111100010111: DATA = 12'b101011001100;
            14'b11_111100011000: DATA = 12'b101011001001;
            14'b11_111100011001: DATA = 12'b101011000110;
            14'b11_111100011010: DATA = 12'b101011000011;
            14'b11_111100011011: DATA = 12'b101011000000;
            14'b11_111100011100: DATA = 12'b101010111101;
            14'b11_111100011101: DATA = 12'b101010111010;
            14'b11_111100011110: DATA = 12'b101010110111;
            14'b11_111100011111: DATA = 12'b101010110100;
            14'b11_111100100000: DATA = 12'b101010110001;
            14'b11_111100100001: DATA = 12'b101010101110;
            14'b11_111100100010: DATA = 12'b101010101011;
            14'b11_111100100011: DATA = 12'b101010101000;
            14'b11_111100100100: DATA = 12'b101010100101;
            14'b11_111100100101: DATA = 12'b101010100010;
            14'b11_111100100110: DATA = 12'b101010011111;
            14'b11_111100100111: DATA = 12'b101010011100;
            14'b11_111100101000: DATA = 12'b101010011001;
            14'b11_111100101001: DATA = 12'b101010010110;
            14'b11_111100101010: DATA = 12'b101010010011;
            14'b11_111100101011: DATA = 12'b101010010000;
            14'b11_111100101100: DATA = 12'b101010001110;
            14'b11_111100101101: DATA = 12'b101010001011;
            14'b11_111100101110: DATA = 12'b101010001000;
            14'b11_111100101111: DATA = 12'b101010000101;
            14'b11_111100110000: DATA = 12'b101010000010;
            14'b11_111100110001: DATA = 12'b101001111111;
            14'b11_111100110010: DATA = 12'b101001111100;
            14'b11_111100110011: DATA = 12'b101001111001;
            14'b11_111100110100: DATA = 12'b101001110110;
            14'b11_111100110101: DATA = 12'b101001110011;
            14'b11_111100110110: DATA = 12'b101001110000;
            14'b11_111100110111: DATA = 12'b101001101101;
            14'b11_111100111000: DATA = 12'b101001101010;
            14'b11_111100111001: DATA = 12'b101001100111;
            14'b11_111100111010: DATA = 12'b101001100100;
            14'b11_111100111011: DATA = 12'b101001100001;
            14'b11_111100111100: DATA = 12'b101001011110;
            14'b11_111100111101: DATA = 12'b101001011011;
            14'b11_111100111110: DATA = 12'b101001011000;
            14'b11_111100111111: DATA = 12'b101001010101;
            14'b11_111101000000: DATA = 12'b101001010010;
            14'b11_111101000001: DATA = 12'b101001001111;
            14'b11_111101000010: DATA = 12'b101001001100;
            14'b11_111101000011: DATA = 12'b101001001001;
            14'b11_111101000100: DATA = 12'b101001000110;
            14'b11_111101000101: DATA = 12'b101001000011;
            14'b11_111101000110: DATA = 12'b101001000000;
            14'b11_111101000111: DATA = 12'b101000111101;
            14'b11_111101001000: DATA = 12'b101000111010;
            14'b11_111101001001: DATA = 12'b101000110111;
            14'b11_111101001010: DATA = 12'b101000110100;
            14'b11_111101001011: DATA = 12'b101000110001;
            14'b11_111101001100: DATA = 12'b101000101110;
            14'b11_111101001101: DATA = 12'b101000101011;
            14'b11_111101001110: DATA = 12'b101000101000;
            14'b11_111101001111: DATA = 12'b101000100100;
            14'b11_111101010000: DATA = 12'b101000100001;
            14'b11_111101010001: DATA = 12'b101000011110;
            14'b11_111101010010: DATA = 12'b101000011011;
            14'b11_111101010011: DATA = 12'b101000011000;
            14'b11_111101010100: DATA = 12'b101000010101;
            14'b11_111101010101: DATA = 12'b101000010010;
            14'b11_111101010110: DATA = 12'b101000001111;
            14'b11_111101010111: DATA = 12'b101000001100;
            14'b11_111101011000: DATA = 12'b101000001001;
            14'b11_111101011001: DATA = 12'b101000000110;
            14'b11_111101011010: DATA = 12'b101000000011;
            14'b11_111101011011: DATA = 12'b101000000000;
            14'b11_111101011100: DATA = 12'b100111111101;
            14'b11_111101011101: DATA = 12'b100111111010;
            14'b11_111101011110: DATA = 12'b100111110111;
            14'b11_111101011111: DATA = 12'b100111110100;
            14'b11_111101100000: DATA = 12'b100111110001;
            14'b11_111101100001: DATA = 12'b100111101110;
            14'b11_111101100010: DATA = 12'b100111101011;
            14'b11_111101100011: DATA = 12'b100111101000;
            14'b11_111101100100: DATA = 12'b100111100101;
            14'b11_111101100101: DATA = 12'b100111100010;
            14'b11_111101100110: DATA = 12'b100111011111;
            14'b11_111101100111: DATA = 12'b100111011100;
            14'b11_111101101000: DATA = 12'b100111011000;
            14'b11_111101101001: DATA = 12'b100111010101;
            14'b11_111101101010: DATA = 12'b100111010010;
            14'b11_111101101011: DATA = 12'b100111001111;
            14'b11_111101101100: DATA = 12'b100111001100;
            14'b11_111101101101: DATA = 12'b100111001001;
            14'b11_111101101110: DATA = 12'b100111000110;
            14'b11_111101101111: DATA = 12'b100111000011;
            14'b11_111101110000: DATA = 12'b100111000000;
            14'b11_111101110001: DATA = 12'b100110111101;
            14'b11_111101110010: DATA = 12'b100110111010;
            14'b11_111101110011: DATA = 12'b100110110111;
            14'b11_111101110100: DATA = 12'b100110110100;
            14'b11_111101110101: DATA = 12'b100110110001;
            14'b11_111101110110: DATA = 12'b100110101110;
            14'b11_111101110111: DATA = 12'b100110101011;
            14'b11_111101111000: DATA = 12'b100110100111;
            14'b11_111101111001: DATA = 12'b100110100100;
            14'b11_111101111010: DATA = 12'b100110100001;
            14'b11_111101111011: DATA = 12'b100110011110;
            14'b11_111101111100: DATA = 12'b100110011011;
            14'b11_111101111101: DATA = 12'b100110011000;
            14'b11_111101111110: DATA = 12'b100110010101;
            14'b11_111101111111: DATA = 12'b100110010010;
            14'b11_111110000000: DATA = 12'b100110001111;
            14'b11_111110000001: DATA = 12'b100110001100;
            14'b11_111110000010: DATA = 12'b100110001001;
            14'b11_111110000011: DATA = 12'b100110000110;
            14'b11_111110000100: DATA = 12'b100110000011;
            14'b11_111110000101: DATA = 12'b100101111111;
            14'b11_111110000110: DATA = 12'b100101111100;
            14'b11_111110000111: DATA = 12'b100101111001;
            14'b11_111110001000: DATA = 12'b100101110110;
            14'b11_111110001001: DATA = 12'b100101110011;
            14'b11_111110001010: DATA = 12'b100101110000;
            14'b11_111110001011: DATA = 12'b100101101101;
            14'b11_111110001100: DATA = 12'b100101101010;
            14'b11_111110001101: DATA = 12'b100101100111;
            14'b11_111110001110: DATA = 12'b100101100100;
            14'b11_111110001111: DATA = 12'b100101100001;
            14'b11_111110010000: DATA = 12'b100101011101;
            14'b11_111110010001: DATA = 12'b100101011010;
            14'b11_111110010010: DATA = 12'b100101010111;
            14'b11_111110010011: DATA = 12'b100101010100;
            14'b11_111110010100: DATA = 12'b100101010001;
            14'b11_111110010101: DATA = 12'b100101001110;
            14'b11_111110010110: DATA = 12'b100101001011;
            14'b11_111110010111: DATA = 12'b100101001000;
            14'b11_111110011000: DATA = 12'b100101000101;
            14'b11_111110011001: DATA = 12'b100101000010;
            14'b11_111110011010: DATA = 12'b100100111110;
            14'b11_111110011011: DATA = 12'b100100111011;
            14'b11_111110011100: DATA = 12'b100100111000;
            14'b11_111110011101: DATA = 12'b100100110101;
            14'b11_111110011110: DATA = 12'b100100110010;
            14'b11_111110011111: DATA = 12'b100100101111;
            14'b11_111110100000: DATA = 12'b100100101100;
            14'b11_111110100001: DATA = 12'b100100101001;
            14'b11_111110100010: DATA = 12'b100100100110;
            14'b11_111110100011: DATA = 12'b100100100011;
            14'b11_111110100100: DATA = 12'b100100011111;
            14'b11_111110100101: DATA = 12'b100100011100;
            14'b11_111110100110: DATA = 12'b100100011001;
            14'b11_111110100111: DATA = 12'b100100010110;
            14'b11_111110101000: DATA = 12'b100100010011;
            14'b11_111110101001: DATA = 12'b100100010000;
            14'b11_111110101010: DATA = 12'b100100001101;
            14'b11_111110101011: DATA = 12'b100100001010;
            14'b11_111110101100: DATA = 12'b100100000111;
            14'b11_111110101101: DATA = 12'b100100000011;
            14'b11_111110101110: DATA = 12'b100100000000;
            14'b11_111110101111: DATA = 12'b100011111101;
            14'b11_111110110000: DATA = 12'b100011111010;
            14'b11_111110110001: DATA = 12'b100011110111;
            14'b11_111110110010: DATA = 12'b100011110100;
            14'b11_111110110011: DATA = 12'b100011110001;
            14'b11_111110110100: DATA = 12'b100011101110;
            14'b11_111110110101: DATA = 12'b100011101010;
            14'b11_111110110110: DATA = 12'b100011100111;
            14'b11_111110110111: DATA = 12'b100011100100;
            14'b11_111110111000: DATA = 12'b100011100001;
            14'b11_111110111001: DATA = 12'b100011011110;
            14'b11_111110111010: DATA = 12'b100011011011;
            14'b11_111110111011: DATA = 12'b100011011000;
            14'b11_111110111100: DATA = 12'b100011010101;
            14'b11_111110111101: DATA = 12'b100011010010;
            14'b11_111110111110: DATA = 12'b100011001110;
            14'b11_111110111111: DATA = 12'b100011001011;
            14'b11_111111000000: DATA = 12'b100011001000;
            14'b11_111111000001: DATA = 12'b100011000101;
            14'b11_111111000010: DATA = 12'b100011000010;
            14'b11_111111000011: DATA = 12'b100010111111;
            14'b11_111111000100: DATA = 12'b100010111100;
            14'b11_111111000101: DATA = 12'b100010111001;
            14'b11_111111000110: DATA = 12'b100010110101;
            14'b11_111111000111: DATA = 12'b100010110010;
            14'b11_111111001000: DATA = 12'b100010101111;
            14'b11_111111001001: DATA = 12'b100010101100;
            14'b11_111111001010: DATA = 12'b100010101001;
            14'b11_111111001011: DATA = 12'b100010100110;
            14'b11_111111001100: DATA = 12'b100010100011;
            14'b11_111111001101: DATA = 12'b100010011111;
            14'b11_111111001110: DATA = 12'b100010011100;
            14'b11_111111001111: DATA = 12'b100010011001;
            14'b11_111111010000: DATA = 12'b100010010110;
            14'b11_111111010001: DATA = 12'b100010010011;
            14'b11_111111010010: DATA = 12'b100010010000;
            14'b11_111111010011: DATA = 12'b100010001101;
            14'b11_111111010100: DATA = 12'b100010001010;
            14'b11_111111010101: DATA = 12'b100010000110;
            14'b11_111111010110: DATA = 12'b100010000011;
            14'b11_111111010111: DATA = 12'b100010000000;
            14'b11_111111011000: DATA = 12'b100001111101;
            14'b11_111111011001: DATA = 12'b100001111010;
            14'b11_111111011010: DATA = 12'b100001110111;
            14'b11_111111011011: DATA = 12'b100001110100;
            14'b11_111111011100: DATA = 12'b100001110000;
            14'b11_111111011101: DATA = 12'b100001101101;
            14'b11_111111011110: DATA = 12'b100001101010;
            14'b11_111111011111: DATA = 12'b100001100111;
            14'b11_111111100000: DATA = 12'b100001100100;
            14'b11_111111100001: DATA = 12'b100001100001;
            14'b11_111111100010: DATA = 12'b100001011110;
            14'b11_111111100011: DATA = 12'b100001011011;
            14'b11_111111100100: DATA = 12'b100001010111;
            14'b11_111111100101: DATA = 12'b100001010100;
            14'b11_111111100110: DATA = 12'b100001010001;
            14'b11_111111100111: DATA = 12'b100001001110;
            14'b11_111111101000: DATA = 12'b100001001011;
            14'b11_111111101001: DATA = 12'b100001001000;
            14'b11_111111101010: DATA = 12'b100001000101;
            14'b11_111111101011: DATA = 12'b100001000001;
            14'b11_111111101100: DATA = 12'b100000111110;
            14'b11_111111101101: DATA = 12'b100000111011;
            14'b11_111111101110: DATA = 12'b100000111000;
            14'b11_111111101111: DATA = 12'b100000110101;
            14'b11_111111110000: DATA = 12'b100000110010;
            14'b11_111111110001: DATA = 12'b100000101111;
            14'b11_111111110010: DATA = 12'b100000101011;
            14'b11_111111110011: DATA = 12'b100000101000;
            14'b11_111111110100: DATA = 12'b100000100101;
            14'b11_111111110101: DATA = 12'b100000100010;
            14'b11_111111110110: DATA = 12'b100000011111;
            14'b11_111111110111: DATA = 12'b100000011100;
            14'b11_111111111000: DATA = 12'b100000011001;
            14'b11_111111111001: DATA = 12'b100000010101;
            14'b11_111111111010: DATA = 12'b100000010010;
            14'b11_111111111011: DATA = 12'b100000001111;
            14'b11_111111111100: DATA = 12'b100000001100;
            14'b11_111111111101: DATA = 12'b100000001001;
            14'b11_111111111110: DATA = 12'b100000000110;
            14'b11_111111111111: DATA = 12'b100000000011;
        endcase
    end    
endmodule
