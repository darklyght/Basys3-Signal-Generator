`timescale 1ns / 1ps

module bcd_to_ascii_amp(
    input [15:0] BCD,
    output [31:0] ASCII
    );
    
    assign ASCII[7:0] = (BCD[3:0] == 4'b0000) ? 8'h30 :
                            (BCD[3:0] == 4'b0001) ? 8'h31 :
                            (BCD[3:0] == 4'b0010) ? 8'h32 :
                            (BCD[3:0] == 4'b0011) ? 8'h33 :
                            (BCD[3:0] == 4'b0100) ? 8'h34 :
                            (BCD[3:0] == 4'b0101) ? 8'h35 :
                            (BCD[3:0] == 4'b0110) ? 8'h36 :
                            (BCD[3:0] == 4'b0111) ? 8'h37 :
                            (BCD[3:0] == 4'b1000) ? 8'h38 :
                            (BCD[3:0] == 4'b1001) ? 8'h39 : 8'h00;
    assign ASCII[15:8] = (BCD[7:4] == 4'b0000) ? 8'h30 :
                         (BCD[7:4] == 4'b0001) ? 8'h31 :
                         (BCD[7:4] == 4'b0010) ? 8'h32 :
                         (BCD[7:4] == 4'b0011) ? 8'h33 :
                         (BCD[7:4] == 4'b0100) ? 8'h34 :
                         (BCD[7:4] == 4'b0101) ? 8'h35 :
                         (BCD[7:4] == 4'b0110) ? 8'h36 :
                         (BCD[7:4] == 4'b0111) ? 8'h37 :
                         (BCD[7:4] == 4'b1000) ? 8'h38 :
                         (BCD[7:4] == 4'b1001) ? 8'h39 : 8'h00;
    assign ASCII[23:16] = (BCD[11:8] == 4'b0000) ? 8'h30 :
                          (BCD[11:8] == 4'b0001) ? 8'h31 :
                          (BCD[11:8] == 4'b0010) ? 8'h32 :
                          (BCD[11:8] == 4'b0011) ? 8'h33 :
                          (BCD[11:8] == 4'b0100) ? 8'h34 :
                          (BCD[11:8] == 4'b0101) ? 8'h35 :
                          (BCD[11:8] == 4'b0110) ? 8'h36 :
                          (BCD[11:8] == 4'b0111) ? 8'h37 :
                          (BCD[11:8] == 4'b1000) ? 8'h38 :
                          (BCD[11:8] == 4'b1001) ? 8'h39 : 8'h00;
    assign ASCII[31:24] = (BCD[15:12] == 4'b0000) ? 8'h30 :
                          (BCD[15:12] == 4'b0001) ? 8'h31 :
                          (BCD[15:12] == 4'b0010) ? 8'h32 :
                          (BCD[15:12] == 4'b0011) ? 8'h33 :
                          (BCD[15:12] == 4'b0100) ? 8'h34 :
                          (BCD[15:12] == 4'b0101) ? 8'h35 :
                          (BCD[15:12] == 4'b0110) ? 8'h36 :
                          (BCD[15:12] == 4'b0111) ? 8'h37 :
                          (BCD[15:12] == 4'b1000) ? 8'h38 :
                          (BCD[15:12] == 4'b1001) ? 8'h39 : 8'h00;
endmodule
